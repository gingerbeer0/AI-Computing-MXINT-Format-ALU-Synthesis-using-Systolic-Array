`timescale 1ns/1ps

module TOP_tb;
    parameter integer NUM_INPUTS = 256;
    parameter integer NUM_OUTPUTS = 896;
    parameter integer DECIMAL_N0 = 10; // MXINT fixed-point decimal location
    parameter integer DECIMAL_N1 = 8; // Final Result fixed-point decimal location

    logic CLK;
    logic RSTN;
    logic [1:0] calc;
    logic [15:0] inputs[0:NUM_INPUTS-1];
    logic [15:0] MXINT_outputs[0:NUM_INPUTS-1];
    logic [15:0] RESULT_outputs[0:NUM_OUTPUTS-1];

    //logic [15:0] FP16_inputs[0:NUM_INPUTS-1];
    logic [15:0] FP16_expected[0:NUM_OUTPUTS-1];
    real mxint_snr, snr_mult, snr_add, snr_sub;
 
    integer cycle_count_mult, cycle_count_add, cycle_count_sub, cycle_count_mxint;
    integer log_file;

    TOP dut (
        .CLK(CLK),
        .RSTN(RSTN),
        .calc(calc),

        .INPUT_0(inputs[0]),
        .INPUT_1(inputs[1]),
        .INPUT_2(inputs[2]),
        .INPUT_3(inputs[3]),
        .INPUT_4(inputs[4]),
        .INPUT_5(inputs[5]),
        .INPUT_6(inputs[6]),
        .INPUT_7(inputs[7]),
        .INPUT_8(inputs[8]),
        .INPUT_9(inputs[9]),
        .INPUT_10(inputs[10]),
        .INPUT_11(inputs[11]),
        .INPUT_12(inputs[12]),
        .INPUT_13(inputs[13]),
        .INPUT_14(inputs[14]),
        .INPUT_15(inputs[15]),
        .INPUT_16(inputs[16]),
        .INPUT_17(inputs[17]),
        .INPUT_18(inputs[18]),
        .INPUT_19(inputs[19]),
        .INPUT_20(inputs[20]),
        .INPUT_21(inputs[21]),
        .INPUT_22(inputs[22]),
        .INPUT_23(inputs[23]),
        .INPUT_24(inputs[24]),
        .INPUT_25(inputs[25]),
        .INPUT_26(inputs[26]),
        .INPUT_27(inputs[27]),
        .INPUT_28(inputs[28]),
        .INPUT_29(inputs[29]),
        .INPUT_30(inputs[30]),
        .INPUT_31(inputs[31]),
        .INPUT_32(inputs[32]),
        .INPUT_33(inputs[33]),
        .INPUT_34(inputs[34]),
        .INPUT_35(inputs[35]),
        .INPUT_36(inputs[36]),
        .INPUT_37(inputs[37]),
        .INPUT_38(inputs[38]),
        .INPUT_39(inputs[39]),
        .INPUT_40(inputs[40]),
        .INPUT_41(inputs[41]),
        .INPUT_42(inputs[42]),
        .INPUT_43(inputs[43]),
        .INPUT_44(inputs[44]),
        .INPUT_45(inputs[45]),
        .INPUT_46(inputs[46]),
        .INPUT_47(inputs[47]),
        .INPUT_48(inputs[48]),
        .INPUT_49(inputs[49]),
        .INPUT_50(inputs[50]),
        .INPUT_51(inputs[51]),
        .INPUT_52(inputs[52]),
        .INPUT_53(inputs[53]),
        .INPUT_54(inputs[54]),
        .INPUT_55(inputs[55]),
        .INPUT_56(inputs[56]),
        .INPUT_57(inputs[57]),
        .INPUT_58(inputs[58]),
        .INPUT_59(inputs[59]),
        .INPUT_60(inputs[60]),
        .INPUT_61(inputs[61]),
        .INPUT_62(inputs[62]),
        .INPUT_63(inputs[63]),
        .INPUT_64(inputs[64]),
        .INPUT_65(inputs[65]),
        .INPUT_66(inputs[66]),
        .INPUT_67(inputs[67]),
        .INPUT_68(inputs[68]),
        .INPUT_69(inputs[69]),
        .INPUT_70(inputs[70]),
        .INPUT_71(inputs[71]),
        .INPUT_72(inputs[72]),
        .INPUT_73(inputs[73]),
        .INPUT_74(inputs[74]),
        .INPUT_75(inputs[75]),
        .INPUT_76(inputs[76]),
        .INPUT_77(inputs[77]),
        .INPUT_78(inputs[78]),
        .INPUT_79(inputs[79]),
        .INPUT_80(inputs[80]),
        .INPUT_81(inputs[81]),
        .INPUT_82(inputs[82]),
        .INPUT_83(inputs[83]),
        .INPUT_84(inputs[84]),
        .INPUT_85(inputs[85]),
        .INPUT_86(inputs[86]),
        .INPUT_87(inputs[87]),
        .INPUT_88(inputs[88]),
        .INPUT_89(inputs[89]),
        .INPUT_90(inputs[90]),
        .INPUT_91(inputs[91]),
        .INPUT_92(inputs[92]),
        .INPUT_93(inputs[93]),
        .INPUT_94(inputs[94]),
        .INPUT_95(inputs[95]),
        .INPUT_96(inputs[96]),
        .INPUT_97(inputs[97]),
        .INPUT_98(inputs[98]),
        .INPUT_99(inputs[99]),
        .INPUT_100(inputs[100]),
        .INPUT_101(inputs[101]),
        .INPUT_102(inputs[102]),
        .INPUT_103(inputs[103]),
        .INPUT_104(inputs[104]),
        .INPUT_105(inputs[105]),
        .INPUT_106(inputs[106]),
        .INPUT_107(inputs[107]),
        .INPUT_108(inputs[108]),
        .INPUT_109(inputs[109]),
        .INPUT_110(inputs[110]),
        .INPUT_111(inputs[111]),
        .INPUT_112(inputs[112]),
        .INPUT_113(inputs[113]),
        .INPUT_114(inputs[114]),
        .INPUT_115(inputs[115]),
        .INPUT_116(inputs[116]),
        .INPUT_117(inputs[117]),
        .INPUT_118(inputs[118]),
        .INPUT_119(inputs[119]),
        .INPUT_120(inputs[120]),
        .INPUT_121(inputs[121]),
        .INPUT_122(inputs[122]),
        .INPUT_123(inputs[123]),
        .INPUT_124(inputs[124]),
        .INPUT_125(inputs[125]),
        .INPUT_126(inputs[126]),
        .INPUT_127(inputs[127]),
        .INPUT_128(inputs[128]),
        .INPUT_129(inputs[129]),
        .INPUT_130(inputs[130]),
        .INPUT_131(inputs[131]),
        .INPUT_132(inputs[132]),
        .INPUT_133(inputs[133]),
        .INPUT_134(inputs[134]),
        .INPUT_135(inputs[135]),
        .INPUT_136(inputs[136]),
        .INPUT_137(inputs[137]),
        .INPUT_138(inputs[138]),
        .INPUT_139(inputs[139]),
        .INPUT_140(inputs[140]),
        .INPUT_141(inputs[141]),
        .INPUT_142(inputs[142]),
        .INPUT_143(inputs[143]),
        .INPUT_144(inputs[144]),
        .INPUT_145(inputs[145]),
        .INPUT_146(inputs[146]),
        .INPUT_147(inputs[147]),
        .INPUT_148(inputs[148]),
        .INPUT_149(inputs[149]),
        .INPUT_150(inputs[150]),
        .INPUT_151(inputs[151]),
        .INPUT_152(inputs[152]),
        .INPUT_153(inputs[153]),
        .INPUT_154(inputs[154]),
        .INPUT_155(inputs[155]),
        .INPUT_156(inputs[156]),
        .INPUT_157(inputs[157]),
        .INPUT_158(inputs[158]),
        .INPUT_159(inputs[159]),
        .INPUT_160(inputs[160]),
        .INPUT_161(inputs[161]),
        .INPUT_162(inputs[162]),
        .INPUT_163(inputs[163]),
        .INPUT_164(inputs[164]),
        .INPUT_165(inputs[165]),
        .INPUT_166(inputs[166]),
        .INPUT_167(inputs[167]),
        .INPUT_168(inputs[168]),
        .INPUT_169(inputs[169]),
        .INPUT_170(inputs[170]),
        .INPUT_171(inputs[171]),
        .INPUT_172(inputs[172]),
        .INPUT_173(inputs[173]),
        .INPUT_174(inputs[174]),
        .INPUT_175(inputs[175]),
        .INPUT_176(inputs[176]),
        .INPUT_177(inputs[177]),
        .INPUT_178(inputs[178]),
        .INPUT_179(inputs[179]),
        .INPUT_180(inputs[180]),
        .INPUT_181(inputs[181]),
        .INPUT_182(inputs[182]),
        .INPUT_183(inputs[183]),
        .INPUT_184(inputs[184]),
        .INPUT_185(inputs[185]),
        .INPUT_186(inputs[186]),
        .INPUT_187(inputs[187]),
        .INPUT_188(inputs[188]),
        .INPUT_189(inputs[189]),
        .INPUT_190(inputs[190]),
        .INPUT_191(inputs[191]),
        .INPUT_192(inputs[192]),
        .INPUT_193(inputs[193]),
        .INPUT_194(inputs[194]),
        .INPUT_195(inputs[195]),
        .INPUT_196(inputs[196]),
        .INPUT_197(inputs[197]),
        .INPUT_198(inputs[198]),
        .INPUT_199(inputs[199]),
        .INPUT_200(inputs[200]),
        .INPUT_201(inputs[201]),
        .INPUT_202(inputs[202]),
        .INPUT_203(inputs[203]),
        .INPUT_204(inputs[204]),
        .INPUT_205(inputs[205]),
        .INPUT_206(inputs[206]),
        .INPUT_207(inputs[207]),
        .INPUT_208(inputs[208]),
        .INPUT_209(inputs[209]),
        .INPUT_210(inputs[210]),
        .INPUT_211(inputs[211]),
        .INPUT_212(inputs[212]),
        .INPUT_213(inputs[213]),
        .INPUT_214(inputs[214]),
        .INPUT_215(inputs[215]),
        .INPUT_216(inputs[216]),
        .INPUT_217(inputs[217]),
        .INPUT_218(inputs[218]),
        .INPUT_219(inputs[219]),
        .INPUT_220(inputs[220]),
        .INPUT_221(inputs[221]),
        .INPUT_222(inputs[222]),
        .INPUT_223(inputs[223]),
        .INPUT_224(inputs[224]),
        .INPUT_225(inputs[225]),
        .INPUT_226(inputs[226]),
        .INPUT_227(inputs[227]),
        .INPUT_228(inputs[228]),
        .INPUT_229(inputs[229]),
        .INPUT_230(inputs[230]),
        .INPUT_231(inputs[231]),
        .INPUT_232(inputs[232]),
        .INPUT_233(inputs[233]),
        .INPUT_234(inputs[234]),
        .INPUT_235(inputs[235]),
        .INPUT_236(inputs[236]),
        .INPUT_237(inputs[237]),
        .INPUT_238(inputs[238]),
        .INPUT_239(inputs[239]),
        .INPUT_240(inputs[240]),
        .INPUT_241(inputs[241]),
        .INPUT_242(inputs[242]),
        .INPUT_243(inputs[243]),
        .INPUT_244(inputs[244]),
        .INPUT_245(inputs[245]),
        .INPUT_246(inputs[246]),
        .INPUT_247(inputs[247]),
        .INPUT_248(inputs[248]),
        .INPUT_249(inputs[249]),
        .INPUT_250(inputs[250]),
        .INPUT_251(inputs[251]),
        .INPUT_252(inputs[252]),
        .INPUT_253(inputs[253]),
        .INPUT_254(inputs[254]),
        .INPUT_255(inputs[255]),


        .MXINT_0(MXINT_outputs[0]),
        .MXINT_1(MXINT_outputs[1]),
        .MXINT_2(MXINT_outputs[2]),
        .MXINT_3(MXINT_outputs[3]),
        .MXINT_4(MXINT_outputs[4]),
        .MXINT_5(MXINT_outputs[5]),
        .MXINT_6(MXINT_outputs[6]),
        .MXINT_7(MXINT_outputs[7]),
        .MXINT_8(MXINT_outputs[8]),
        .MXINT_9(MXINT_outputs[9]),
        .MXINT_10(MXINT_outputs[10]),
        .MXINT_11(MXINT_outputs[11]),
        .MXINT_12(MXINT_outputs[12]),
        .MXINT_13(MXINT_outputs[13]),
        .MXINT_14(MXINT_outputs[14]),
        .MXINT_15(MXINT_outputs[15]),
        .MXINT_16(MXINT_outputs[16]),
        .MXINT_17(MXINT_outputs[17]),
        .MXINT_18(MXINT_outputs[18]),
        .MXINT_19(MXINT_outputs[19]),
        .MXINT_20(MXINT_outputs[20]),
        .MXINT_21(MXINT_outputs[21]),
        .MXINT_22(MXINT_outputs[22]),
        .MXINT_23(MXINT_outputs[23]),
        .MXINT_24(MXINT_outputs[24]),
        .MXINT_25(MXINT_outputs[25]),
        .MXINT_26(MXINT_outputs[26]),
        .MXINT_27(MXINT_outputs[27]),
        .MXINT_28(MXINT_outputs[28]),
        .MXINT_29(MXINT_outputs[29]),
        .MXINT_30(MXINT_outputs[30]),
        .MXINT_31(MXINT_outputs[31]),
        .MXINT_32(MXINT_outputs[32]),
        .MXINT_33(MXINT_outputs[33]),
        .MXINT_34(MXINT_outputs[34]),
        .MXINT_35(MXINT_outputs[35]),
        .MXINT_36(MXINT_outputs[36]),
        .MXINT_37(MXINT_outputs[37]),
        .MXINT_38(MXINT_outputs[38]),
        .MXINT_39(MXINT_outputs[39]),
        .MXINT_40(MXINT_outputs[40]),
        .MXINT_41(MXINT_outputs[41]),
        .MXINT_42(MXINT_outputs[42]),
        .MXINT_43(MXINT_outputs[43]),
        .MXINT_44(MXINT_outputs[44]),
        .MXINT_45(MXINT_outputs[45]),
        .MXINT_46(MXINT_outputs[46]),
        .MXINT_47(MXINT_outputs[47]),
        .MXINT_48(MXINT_outputs[48]),
        .MXINT_49(MXINT_outputs[49]),
        .MXINT_50(MXINT_outputs[50]),
        .MXINT_51(MXINT_outputs[51]),
        .MXINT_52(MXINT_outputs[52]),
        .MXINT_53(MXINT_outputs[53]),
        .MXINT_54(MXINT_outputs[54]),
        .MXINT_55(MXINT_outputs[55]),
        .MXINT_56(MXINT_outputs[56]),
        .MXINT_57(MXINT_outputs[57]),
        .MXINT_58(MXINT_outputs[58]),
        .MXINT_59(MXINT_outputs[59]),
        .MXINT_60(MXINT_outputs[60]),
        .MXINT_61(MXINT_outputs[61]),
        .MXINT_62(MXINT_outputs[62]),
        .MXINT_63(MXINT_outputs[63]),
        .MXINT_64(MXINT_outputs[64]),
        .MXINT_65(MXINT_outputs[65]),
        .MXINT_66(MXINT_outputs[66]),
        .MXINT_67(MXINT_outputs[67]),
        .MXINT_68(MXINT_outputs[68]),
        .MXINT_69(MXINT_outputs[69]),
        .MXINT_70(MXINT_outputs[70]),
        .MXINT_71(MXINT_outputs[71]),
        .MXINT_72(MXINT_outputs[72]),
        .MXINT_73(MXINT_outputs[73]),
        .MXINT_74(MXINT_outputs[74]),
        .MXINT_75(MXINT_outputs[75]),
        .MXINT_76(MXINT_outputs[76]),
        .MXINT_77(MXINT_outputs[77]),
        .MXINT_78(MXINT_outputs[78]),
        .MXINT_79(MXINT_outputs[79]),
        .MXINT_80(MXINT_outputs[80]),
        .MXINT_81(MXINT_outputs[81]),
        .MXINT_82(MXINT_outputs[82]),
        .MXINT_83(MXINT_outputs[83]),
        .MXINT_84(MXINT_outputs[84]),
        .MXINT_85(MXINT_outputs[85]),
        .MXINT_86(MXINT_outputs[86]),
        .MXINT_87(MXINT_outputs[87]),
        .MXINT_88(MXINT_outputs[88]),
        .MXINT_89(MXINT_outputs[89]),
        .MXINT_90(MXINT_outputs[90]),
        .MXINT_91(MXINT_outputs[91]),
        .MXINT_92(MXINT_outputs[92]),
        .MXINT_93(MXINT_outputs[93]),
        .MXINT_94(MXINT_outputs[94]),
        .MXINT_95(MXINT_outputs[95]),
        .MXINT_96(MXINT_outputs[96]),
        .MXINT_97(MXINT_outputs[97]),
        .MXINT_98(MXINT_outputs[98]),
        .MXINT_99(MXINT_outputs[99]),
        .MXINT_100(MXINT_outputs[100]),
        .MXINT_101(MXINT_outputs[101]),
        .MXINT_102(MXINT_outputs[102]),
        .MXINT_103(MXINT_outputs[103]),
        .MXINT_104(MXINT_outputs[104]),
        .MXINT_105(MXINT_outputs[105]),
        .MXINT_106(MXINT_outputs[106]),
        .MXINT_107(MXINT_outputs[107]),
        .MXINT_108(MXINT_outputs[108]),
        .MXINT_109(MXINT_outputs[109]),
        .MXINT_110(MXINT_outputs[110]),
        .MXINT_111(MXINT_outputs[111]),
        .MXINT_112(MXINT_outputs[112]),
        .MXINT_113(MXINT_outputs[113]),
        .MXINT_114(MXINT_outputs[114]),
        .MXINT_115(MXINT_outputs[115]),
        .MXINT_116(MXINT_outputs[116]),
        .MXINT_117(MXINT_outputs[117]),
        .MXINT_118(MXINT_outputs[118]),
        .MXINT_119(MXINT_outputs[119]),
        .MXINT_120(MXINT_outputs[120]),
        .MXINT_121(MXINT_outputs[121]),
        .MXINT_122(MXINT_outputs[122]),
        .MXINT_123(MXINT_outputs[123]),
        .MXINT_124(MXINT_outputs[124]),
        .MXINT_125(MXINT_outputs[125]),
        .MXINT_126(MXINT_outputs[126]),
        .MXINT_127(MXINT_outputs[127]),
        .MXINT_128(MXINT_outputs[128]),
        .MXINT_129(MXINT_outputs[129]),
        .MXINT_130(MXINT_outputs[130]),
        .MXINT_131(MXINT_outputs[131]),
        .MXINT_132(MXINT_outputs[132]),
        .MXINT_133(MXINT_outputs[133]),
        .MXINT_134(MXINT_outputs[134]),
        .MXINT_135(MXINT_outputs[135]),
        .MXINT_136(MXINT_outputs[136]),
        .MXINT_137(MXINT_outputs[137]),
        .MXINT_138(MXINT_outputs[138]),
        .MXINT_139(MXINT_outputs[139]),
        .MXINT_140(MXINT_outputs[140]),
        .MXINT_141(MXINT_outputs[141]),
        .MXINT_142(MXINT_outputs[142]),
        .MXINT_143(MXINT_outputs[143]),
        .MXINT_144(MXINT_outputs[144]),
        .MXINT_145(MXINT_outputs[145]),
        .MXINT_146(MXINT_outputs[146]),
        .MXINT_147(MXINT_outputs[147]),
        .MXINT_148(MXINT_outputs[148]),
        .MXINT_149(MXINT_outputs[149]),
        .MXINT_150(MXINT_outputs[150]),
        .MXINT_151(MXINT_outputs[151]),
        .MXINT_152(MXINT_outputs[152]),
        .MXINT_153(MXINT_outputs[153]),
        .MXINT_154(MXINT_outputs[154]),
        .MXINT_155(MXINT_outputs[155]),
        .MXINT_156(MXINT_outputs[156]),
        .MXINT_157(MXINT_outputs[157]),
        .MXINT_158(MXINT_outputs[158]),
        .MXINT_159(MXINT_outputs[159]),
        .MXINT_160(MXINT_outputs[160]),
        .MXINT_161(MXINT_outputs[161]),
        .MXINT_162(MXINT_outputs[162]),
        .MXINT_163(MXINT_outputs[163]),
        .MXINT_164(MXINT_outputs[164]),
        .MXINT_165(MXINT_outputs[165]),
        .MXINT_166(MXINT_outputs[166]),
        .MXINT_167(MXINT_outputs[167]),
        .MXINT_168(MXINT_outputs[168]),
        .MXINT_169(MXINT_outputs[169]),
        .MXINT_170(MXINT_outputs[170]),
        .MXINT_171(MXINT_outputs[171]),
        .MXINT_172(MXINT_outputs[172]),
        .MXINT_173(MXINT_outputs[173]),
        .MXINT_174(MXINT_outputs[174]),
        .MXINT_175(MXINT_outputs[175]),
        .MXINT_176(MXINT_outputs[176]),
        .MXINT_177(MXINT_outputs[177]),
        .MXINT_178(MXINT_outputs[178]),
        .MXINT_179(MXINT_outputs[179]),
        .MXINT_180(MXINT_outputs[180]),
        .MXINT_181(MXINT_outputs[181]),
        .MXINT_182(MXINT_outputs[182]),
        .MXINT_183(MXINT_outputs[183]),
        .MXINT_184(MXINT_outputs[184]),
        .MXINT_185(MXINT_outputs[185]),
        .MXINT_186(MXINT_outputs[186]),
        .MXINT_187(MXINT_outputs[187]),
        .MXINT_188(MXINT_outputs[188]),
        .MXINT_189(MXINT_outputs[189]),
        .MXINT_190(MXINT_outputs[190]),
        .MXINT_191(MXINT_outputs[191]),
        .MXINT_192(MXINT_outputs[192]),
        .MXINT_193(MXINT_outputs[193]),
        .MXINT_194(MXINT_outputs[194]),
        .MXINT_195(MXINT_outputs[195]),
        .MXINT_196(MXINT_outputs[196]),
        .MXINT_197(MXINT_outputs[197]),
        .MXINT_198(MXINT_outputs[198]),
        .MXINT_199(MXINT_outputs[199]),
        .MXINT_200(MXINT_outputs[200]),
        .MXINT_201(MXINT_outputs[201]),
        .MXINT_202(MXINT_outputs[202]),
        .MXINT_203(MXINT_outputs[203]),
        .MXINT_204(MXINT_outputs[204]),
        .MXINT_205(MXINT_outputs[205]),
        .MXINT_206(MXINT_outputs[206]),
        .MXINT_207(MXINT_outputs[207]),
        .MXINT_208(MXINT_outputs[208]),
        .MXINT_209(MXINT_outputs[209]),
        .MXINT_210(MXINT_outputs[210]),
        .MXINT_211(MXINT_outputs[211]),
        .MXINT_212(MXINT_outputs[212]),
        .MXINT_213(MXINT_outputs[213]),
        .MXINT_214(MXINT_outputs[214]),
        .MXINT_215(MXINT_outputs[215]),
        .MXINT_216(MXINT_outputs[216]),
        .MXINT_217(MXINT_outputs[217]),
        .MXINT_218(MXINT_outputs[218]),
        .MXINT_219(MXINT_outputs[219]),
        .MXINT_220(MXINT_outputs[220]),
        .MXINT_221(MXINT_outputs[221]),
        .MXINT_222(MXINT_outputs[222]),
        .MXINT_223(MXINT_outputs[223]),
        .MXINT_224(MXINT_outputs[224]),
        .MXINT_225(MXINT_outputs[225]),
        .MXINT_226(MXINT_outputs[226]),
        .MXINT_227(MXINT_outputs[227]),
        .MXINT_228(MXINT_outputs[228]),
        .MXINT_229(MXINT_outputs[229]),
        .MXINT_230(MXINT_outputs[230]),
        .MXINT_231(MXINT_outputs[231]),
        .MXINT_232(MXINT_outputs[232]),
        .MXINT_233(MXINT_outputs[233]),
        .MXINT_234(MXINT_outputs[234]),
        .MXINT_235(MXINT_outputs[235]),
        .MXINT_236(MXINT_outputs[236]),
        .MXINT_237(MXINT_outputs[237]),
        .MXINT_238(MXINT_outputs[238]),
        .MXINT_239(MXINT_outputs[239]),
        .MXINT_240(MXINT_outputs[240]),
        .MXINT_241(MXINT_outputs[241]),
        .MXINT_242(MXINT_outputs[242]),
        .MXINT_243(MXINT_outputs[243]),
        .MXINT_244(MXINT_outputs[244]),
        .MXINT_245(MXINT_outputs[245]),
        .MXINT_246(MXINT_outputs[246]),
        .MXINT_247(MXINT_outputs[247]),
        .MXINT_248(MXINT_outputs[248]),
        .MXINT_249(MXINT_outputs[249]),
        .MXINT_250(MXINT_outputs[250]),
        .MXINT_251(MXINT_outputs[251]),
        .MXINT_252(MXINT_outputs[252]),
        .MXINT_253(MXINT_outputs[253]),
        .MXINT_254(MXINT_outputs[254]),
        .MXINT_255(MXINT_outputs[255]),


        .RESULT_0(RESULT_outputs[0]),
        .RESULT_1(RESULT_outputs[1]),
        .RESULT_2(RESULT_outputs[2]),
        .RESULT_3(RESULT_outputs[3]),
        .RESULT_4(RESULT_outputs[4]),
        .RESULT_5(RESULT_outputs[5]),
        .RESULT_6(RESULT_outputs[6]),
        .RESULT_7(RESULT_outputs[7]),
        .RESULT_8(RESULT_outputs[8]),
        .RESULT_9(RESULT_outputs[9]),
        .RESULT_10(RESULT_outputs[10]),
        .RESULT_11(RESULT_outputs[11]),
        .RESULT_12(RESULT_outputs[12]),
        .RESULT_13(RESULT_outputs[13]),
        .RESULT_14(RESULT_outputs[14]),
        .RESULT_15(RESULT_outputs[15]),
        .RESULT_16(RESULT_outputs[16]),
        .RESULT_17(RESULT_outputs[17]),
        .RESULT_18(RESULT_outputs[18]),
        .RESULT_19(RESULT_outputs[19]),
        .RESULT_20(RESULT_outputs[20]),
        .RESULT_21(RESULT_outputs[21]),
        .RESULT_22(RESULT_outputs[22]),
        .RESULT_23(RESULT_outputs[23]),
        .RESULT_24(RESULT_outputs[24]),
        .RESULT_25(RESULT_outputs[25]),
        .RESULT_26(RESULT_outputs[26]),
        .RESULT_27(RESULT_outputs[27]),
        .RESULT_28(RESULT_outputs[28]),
        .RESULT_29(RESULT_outputs[29]),
        .RESULT_30(RESULT_outputs[30]),
        .RESULT_31(RESULT_outputs[31]),
        .RESULT_32(RESULT_outputs[32]),
        .RESULT_33(RESULT_outputs[33]),
        .RESULT_34(RESULT_outputs[34]),
        .RESULT_35(RESULT_outputs[35]),
        .RESULT_36(RESULT_outputs[36]),
        .RESULT_37(RESULT_outputs[37]),
        .RESULT_38(RESULT_outputs[38]),
        .RESULT_39(RESULT_outputs[39]),
        .RESULT_40(RESULT_outputs[40]),
        .RESULT_41(RESULT_outputs[41]),
        .RESULT_42(RESULT_outputs[42]),
        .RESULT_43(RESULT_outputs[43]),
        .RESULT_44(RESULT_outputs[44]),
        .RESULT_45(RESULT_outputs[45]),
        .RESULT_46(RESULT_outputs[46]),
        .RESULT_47(RESULT_outputs[47]),
        .RESULT_48(RESULT_outputs[48]),
        .RESULT_49(RESULT_outputs[49]),
        .RESULT_50(RESULT_outputs[50]),
        .RESULT_51(RESULT_outputs[51]),
        .RESULT_52(RESULT_outputs[52]),
        .RESULT_53(RESULT_outputs[53]),
        .RESULT_54(RESULT_outputs[54]),
        .RESULT_55(RESULT_outputs[55]),
        .RESULT_56(RESULT_outputs[56]),
        .RESULT_57(RESULT_outputs[57]),
        .RESULT_58(RESULT_outputs[58]),
        .RESULT_59(RESULT_outputs[59]),
        .RESULT_60(RESULT_outputs[60]),
        .RESULT_61(RESULT_outputs[61]),
        .RESULT_62(RESULT_outputs[62]),
        .RESULT_63(RESULT_outputs[63]),
        .RESULT_64(RESULT_outputs[64]),
        .RESULT_65(RESULT_outputs[65]),
        .RESULT_66(RESULT_outputs[66]),
        .RESULT_67(RESULT_outputs[67]),
        .RESULT_68(RESULT_outputs[68]),
        .RESULT_69(RESULT_outputs[69]),
        .RESULT_70(RESULT_outputs[70]),
        .RESULT_71(RESULT_outputs[71]),
        .RESULT_72(RESULT_outputs[72]),
        .RESULT_73(RESULT_outputs[73]),
        .RESULT_74(RESULT_outputs[74]),
        .RESULT_75(RESULT_outputs[75]),
        .RESULT_76(RESULT_outputs[76]),
        .RESULT_77(RESULT_outputs[77]),
        .RESULT_78(RESULT_outputs[78]),
        .RESULT_79(RESULT_outputs[79]),
        .RESULT_80(RESULT_outputs[80]),
        .RESULT_81(RESULT_outputs[81]),
        .RESULT_82(RESULT_outputs[82]),
        .RESULT_83(RESULT_outputs[83]),
        .RESULT_84(RESULT_outputs[84]),
        .RESULT_85(RESULT_outputs[85]),
        .RESULT_86(RESULT_outputs[86]),
        .RESULT_87(RESULT_outputs[87]),
        .RESULT_88(RESULT_outputs[88]),
        .RESULT_89(RESULT_outputs[89]),
        .RESULT_90(RESULT_outputs[90]),
        .RESULT_91(RESULT_outputs[91]),
        .RESULT_92(RESULT_outputs[92]),
        .RESULT_93(RESULT_outputs[93]),
        .RESULT_94(RESULT_outputs[94]),
        .RESULT_95(RESULT_outputs[95]),
        .RESULT_96(RESULT_outputs[96]),
        .RESULT_97(RESULT_outputs[97]),
        .RESULT_98(RESULT_outputs[98]),
        .RESULT_99(RESULT_outputs[99]),
        .RESULT_100(RESULT_outputs[100]),
        .RESULT_101(RESULT_outputs[101]),
        .RESULT_102(RESULT_outputs[102]),
        .RESULT_103(RESULT_outputs[103]),
        .RESULT_104(RESULT_outputs[104]),
        .RESULT_105(RESULT_outputs[105]),
        .RESULT_106(RESULT_outputs[106]),
        .RESULT_107(RESULT_outputs[107]),
        .RESULT_108(RESULT_outputs[108]),
        .RESULT_109(RESULT_outputs[109]),
        .RESULT_110(RESULT_outputs[110]),
        .RESULT_111(RESULT_outputs[111]),
        .RESULT_112(RESULT_outputs[112]),
        .RESULT_113(RESULT_outputs[113]),
        .RESULT_114(RESULT_outputs[114]),
        .RESULT_115(RESULT_outputs[115]),
        .RESULT_116(RESULT_outputs[116]),
        .RESULT_117(RESULT_outputs[117]),
        .RESULT_118(RESULT_outputs[118]),
        .RESULT_119(RESULT_outputs[119]),
        .RESULT_120(RESULT_outputs[120]),
        .RESULT_121(RESULT_outputs[121]),
        .RESULT_122(RESULT_outputs[122]),
        .RESULT_123(RESULT_outputs[123]),
        .RESULT_124(RESULT_outputs[124]),
        .RESULT_125(RESULT_outputs[125]),
        .RESULT_126(RESULT_outputs[126]),
        .RESULT_127(RESULT_outputs[127]),
        .RESULT_128(RESULT_outputs[128]),
        .RESULT_129(RESULT_outputs[129]),
        .RESULT_130(RESULT_outputs[130]),
        .RESULT_131(RESULT_outputs[131]),
        .RESULT_132(RESULT_outputs[132]),
        .RESULT_133(RESULT_outputs[133]),
        .RESULT_134(RESULT_outputs[134]),
        .RESULT_135(RESULT_outputs[135]),
        .RESULT_136(RESULT_outputs[136]),
        .RESULT_137(RESULT_outputs[137]),
        .RESULT_138(RESULT_outputs[138]),
        .RESULT_139(RESULT_outputs[139]),
        .RESULT_140(RESULT_outputs[140]),
        .RESULT_141(RESULT_outputs[141]),
        .RESULT_142(RESULT_outputs[142]),
        .RESULT_143(RESULT_outputs[143]),
        .RESULT_144(RESULT_outputs[144]),
        .RESULT_145(RESULT_outputs[145]),
        .RESULT_146(RESULT_outputs[146]),
        .RESULT_147(RESULT_outputs[147]),
        .RESULT_148(RESULT_outputs[148]),
        .RESULT_149(RESULT_outputs[149]),
        .RESULT_150(RESULT_outputs[150]),
        .RESULT_151(RESULT_outputs[151]),
        .RESULT_152(RESULT_outputs[152]),
        .RESULT_153(RESULT_outputs[153]),
        .RESULT_154(RESULT_outputs[154]),
        .RESULT_155(RESULT_outputs[155]),
        .RESULT_156(RESULT_outputs[156]),
        .RESULT_157(RESULT_outputs[157]),
        .RESULT_158(RESULT_outputs[158]),
        .RESULT_159(RESULT_outputs[159]),
        .RESULT_160(RESULT_outputs[160]),
        .RESULT_161(RESULT_outputs[161]),
        .RESULT_162(RESULT_outputs[162]),
        .RESULT_163(RESULT_outputs[163]),
        .RESULT_164(RESULT_outputs[164]),
        .RESULT_165(RESULT_outputs[165]),
        .RESULT_166(RESULT_outputs[166]),
        .RESULT_167(RESULT_outputs[167]),
        .RESULT_168(RESULT_outputs[168]),
        .RESULT_169(RESULT_outputs[169]),
        .RESULT_170(RESULT_outputs[170]),
        .RESULT_171(RESULT_outputs[171]),
        .RESULT_172(RESULT_outputs[172]),
        .RESULT_173(RESULT_outputs[173]),
        .RESULT_174(RESULT_outputs[174]),
        .RESULT_175(RESULT_outputs[175]),
        .RESULT_176(RESULT_outputs[176]),
        .RESULT_177(RESULT_outputs[177]),
        .RESULT_178(RESULT_outputs[178]),
        .RESULT_179(RESULT_outputs[179]),
        .RESULT_180(RESULT_outputs[180]),
        .RESULT_181(RESULT_outputs[181]),
        .RESULT_182(RESULT_outputs[182]),
        .RESULT_183(RESULT_outputs[183]),
        .RESULT_184(RESULT_outputs[184]),
        .RESULT_185(RESULT_outputs[185]),
        .RESULT_186(RESULT_outputs[186]),
        .RESULT_187(RESULT_outputs[187]),
        .RESULT_188(RESULT_outputs[188]),
        .RESULT_189(RESULT_outputs[189]),
        .RESULT_190(RESULT_outputs[190]),
        .RESULT_191(RESULT_outputs[191]),
        .RESULT_192(RESULT_outputs[192]),
        .RESULT_193(RESULT_outputs[193]),
        .RESULT_194(RESULT_outputs[194]),
        .RESULT_195(RESULT_outputs[195]),
        .RESULT_196(RESULT_outputs[196]),
        .RESULT_197(RESULT_outputs[197]),
        .RESULT_198(RESULT_outputs[198]),
        .RESULT_199(RESULT_outputs[199]),
        .RESULT_200(RESULT_outputs[200]),
        .RESULT_201(RESULT_outputs[201]),
        .RESULT_202(RESULT_outputs[202]),
        .RESULT_203(RESULT_outputs[203]),
        .RESULT_204(RESULT_outputs[204]),
        .RESULT_205(RESULT_outputs[205]),
        .RESULT_206(RESULT_outputs[206]),
        .RESULT_207(RESULT_outputs[207]),
        .RESULT_208(RESULT_outputs[208]),
        .RESULT_209(RESULT_outputs[209]),
        .RESULT_210(RESULT_outputs[210]),
        .RESULT_211(RESULT_outputs[211]),
        .RESULT_212(RESULT_outputs[212]),
        .RESULT_213(RESULT_outputs[213]),
        .RESULT_214(RESULT_outputs[214]),
        .RESULT_215(RESULT_outputs[215]),
        .RESULT_216(RESULT_outputs[216]),
        .RESULT_217(RESULT_outputs[217]),
        .RESULT_218(RESULT_outputs[218]),
        .RESULT_219(RESULT_outputs[219]),
        .RESULT_220(RESULT_outputs[220]),
        .RESULT_221(RESULT_outputs[221]),
        .RESULT_222(RESULT_outputs[222]),
        .RESULT_223(RESULT_outputs[223]),
        .RESULT_224(RESULT_outputs[224]),
        .RESULT_225(RESULT_outputs[225]),
        .RESULT_226(RESULT_outputs[226]),
        .RESULT_227(RESULT_outputs[227]),
        .RESULT_228(RESULT_outputs[228]),
        .RESULT_229(RESULT_outputs[229]),
        .RESULT_230(RESULT_outputs[230]),
        .RESULT_231(RESULT_outputs[231]),
        .RESULT_232(RESULT_outputs[232]),
        .RESULT_233(RESULT_outputs[233]),
        .RESULT_234(RESULT_outputs[234]),
        .RESULT_235(RESULT_outputs[235]),
        .RESULT_236(RESULT_outputs[236]),
        .RESULT_237(RESULT_outputs[237]),
        .RESULT_238(RESULT_outputs[238]),
        .RESULT_239(RESULT_outputs[239]),
        .RESULT_240(RESULT_outputs[240]),
        .RESULT_241(RESULT_outputs[241]),
        .RESULT_242(RESULT_outputs[242]),
        .RESULT_243(RESULT_outputs[243]),
        .RESULT_244(RESULT_outputs[244]),
        .RESULT_245(RESULT_outputs[245]),
        .RESULT_246(RESULT_outputs[246]),
        .RESULT_247(RESULT_outputs[247]),
        .RESULT_248(RESULT_outputs[248]),
        .RESULT_249(RESULT_outputs[249]),
        .RESULT_250(RESULT_outputs[250]),
        .RESULT_251(RESULT_outputs[251]),
        .RESULT_252(RESULT_outputs[252]),
        .RESULT_253(RESULT_outputs[253]),
        .RESULT_254(RESULT_outputs[254]),
        .RESULT_255(RESULT_outputs[255]),
        .RESULT_256(RESULT_outputs[256]),
        .RESULT_257(RESULT_outputs[257]),
        .RESULT_258(RESULT_outputs[258]),
        .RESULT_259(RESULT_outputs[259]),
        .RESULT_260(RESULT_outputs[260]),
        .RESULT_261(RESULT_outputs[261]),
        .RESULT_262(RESULT_outputs[262]),
        .RESULT_263(RESULT_outputs[263]),
        .RESULT_264(RESULT_outputs[264]),
        .RESULT_265(RESULT_outputs[265]),
        .RESULT_266(RESULT_outputs[266]),
        .RESULT_267(RESULT_outputs[267]),
        .RESULT_268(RESULT_outputs[268]),
        .RESULT_269(RESULT_outputs[269]),
        .RESULT_270(RESULT_outputs[270]),
        .RESULT_271(RESULT_outputs[271]),
        .RESULT_272(RESULT_outputs[272]),
        .RESULT_273(RESULT_outputs[273]),
        .RESULT_274(RESULT_outputs[274]),
        .RESULT_275(RESULT_outputs[275]),
        .RESULT_276(RESULT_outputs[276]),
        .RESULT_277(RESULT_outputs[277]),
        .RESULT_278(RESULT_outputs[278]),
        .RESULT_279(RESULT_outputs[279]),
        .RESULT_280(RESULT_outputs[280]),
        .RESULT_281(RESULT_outputs[281]),
        .RESULT_282(RESULT_outputs[282]),
        .RESULT_283(RESULT_outputs[283]),
        .RESULT_284(RESULT_outputs[284]),
        .RESULT_285(RESULT_outputs[285]),
        .RESULT_286(RESULT_outputs[286]),
        .RESULT_287(RESULT_outputs[287]),
        .RESULT_288(RESULT_outputs[288]),
        .RESULT_289(RESULT_outputs[289]),
        .RESULT_290(RESULT_outputs[290]),
        .RESULT_291(RESULT_outputs[291]),
        .RESULT_292(RESULT_outputs[292]),
        .RESULT_293(RESULT_outputs[293]),
        .RESULT_294(RESULT_outputs[294]),
        .RESULT_295(RESULT_outputs[295]),
        .RESULT_296(RESULT_outputs[296]),
        .RESULT_297(RESULT_outputs[297]),
        .RESULT_298(RESULT_outputs[298]),
        .RESULT_299(RESULT_outputs[299]),
        .RESULT_300(RESULT_outputs[300]),
        .RESULT_301(RESULT_outputs[301]),
        .RESULT_302(RESULT_outputs[302]),
        .RESULT_303(RESULT_outputs[303]),
        .RESULT_304(RESULT_outputs[304]),
        .RESULT_305(RESULT_outputs[305]),
        .RESULT_306(RESULT_outputs[306]),
        .RESULT_307(RESULT_outputs[307]),
        .RESULT_308(RESULT_outputs[308]),
        .RESULT_309(RESULT_outputs[309]),
        .RESULT_310(RESULT_outputs[310]),
        .RESULT_311(RESULT_outputs[311]),
        .RESULT_312(RESULT_outputs[312]),
        .RESULT_313(RESULT_outputs[313]),
        .RESULT_314(RESULT_outputs[314]),
        .RESULT_315(RESULT_outputs[315]),
        .RESULT_316(RESULT_outputs[316]),
        .RESULT_317(RESULT_outputs[317]),
        .RESULT_318(RESULT_outputs[318]),
        .RESULT_319(RESULT_outputs[319]),
        .RESULT_320(RESULT_outputs[320]),
        .RESULT_321(RESULT_outputs[321]),
        .RESULT_322(RESULT_outputs[322]),
        .RESULT_323(RESULT_outputs[323]),
        .RESULT_324(RESULT_outputs[324]),
        .RESULT_325(RESULT_outputs[325]),
        .RESULT_326(RESULT_outputs[326]),
        .RESULT_327(RESULT_outputs[327]),
        .RESULT_328(RESULT_outputs[328]),
        .RESULT_329(RESULT_outputs[329]),
        .RESULT_330(RESULT_outputs[330]),
        .RESULT_331(RESULT_outputs[331]),
        .RESULT_332(RESULT_outputs[332]),
        .RESULT_333(RESULT_outputs[333]),
        .RESULT_334(RESULT_outputs[334]),
        .RESULT_335(RESULT_outputs[335]),
        .RESULT_336(RESULT_outputs[336]),
        .RESULT_337(RESULT_outputs[337]),
        .RESULT_338(RESULT_outputs[338]),
        .RESULT_339(RESULT_outputs[339]),
        .RESULT_340(RESULT_outputs[340]),
        .RESULT_341(RESULT_outputs[341]),
        .RESULT_342(RESULT_outputs[342]),
        .RESULT_343(RESULT_outputs[343]),
        .RESULT_344(RESULT_outputs[344]),
        .RESULT_345(RESULT_outputs[345]),
        .RESULT_346(RESULT_outputs[346]),
        .RESULT_347(RESULT_outputs[347]),
        .RESULT_348(RESULT_outputs[348]),
        .RESULT_349(RESULT_outputs[349]),
        .RESULT_350(RESULT_outputs[350]),
        .RESULT_351(RESULT_outputs[351]),
        .RESULT_352(RESULT_outputs[352]),
        .RESULT_353(RESULT_outputs[353]),
        .RESULT_354(RESULT_outputs[354]),
        .RESULT_355(RESULT_outputs[355]),
        .RESULT_356(RESULT_outputs[356]),
        .RESULT_357(RESULT_outputs[357]),
        .RESULT_358(RESULT_outputs[358]),
        .RESULT_359(RESULT_outputs[359]),
        .RESULT_360(RESULT_outputs[360]),
        .RESULT_361(RESULT_outputs[361]),
        .RESULT_362(RESULT_outputs[362]),
        .RESULT_363(RESULT_outputs[363]),
        .RESULT_364(RESULT_outputs[364]),
        .RESULT_365(RESULT_outputs[365]),
        .RESULT_366(RESULT_outputs[366]),
        .RESULT_367(RESULT_outputs[367]),
        .RESULT_368(RESULT_outputs[368]),
        .RESULT_369(RESULT_outputs[369]),
        .RESULT_370(RESULT_outputs[370]),
        .RESULT_371(RESULT_outputs[371]),
        .RESULT_372(RESULT_outputs[372]),
        .RESULT_373(RESULT_outputs[373]),
        .RESULT_374(RESULT_outputs[374]),
        .RESULT_375(RESULT_outputs[375]),
        .RESULT_376(RESULT_outputs[376]),
        .RESULT_377(RESULT_outputs[377]),
        .RESULT_378(RESULT_outputs[378]),
        .RESULT_379(RESULT_outputs[379]),
        .RESULT_380(RESULT_outputs[380]),
        .RESULT_381(RESULT_outputs[381]),
        .RESULT_382(RESULT_outputs[382]),
        .RESULT_383(RESULT_outputs[383]),
        .RESULT_384(RESULT_outputs[384]),
        .RESULT_385(RESULT_outputs[385]),
        .RESULT_386(RESULT_outputs[386]),
        .RESULT_387(RESULT_outputs[387]),
        .RESULT_388(RESULT_outputs[388]),
        .RESULT_389(RESULT_outputs[389]),
        .RESULT_390(RESULT_outputs[390]),
        .RESULT_391(RESULT_outputs[391]),
        .RESULT_392(RESULT_outputs[392]),
        .RESULT_393(RESULT_outputs[393]),
        .RESULT_394(RESULT_outputs[394]),
        .RESULT_395(RESULT_outputs[395]),
        .RESULT_396(RESULT_outputs[396]),
        .RESULT_397(RESULT_outputs[397]),
        .RESULT_398(RESULT_outputs[398]),
        .RESULT_399(RESULT_outputs[399]),
        .RESULT_400(RESULT_outputs[400]),
        .RESULT_401(RESULT_outputs[401]),
        .RESULT_402(RESULT_outputs[402]),
        .RESULT_403(RESULT_outputs[403]),
        .RESULT_404(RESULT_outputs[404]),
        .RESULT_405(RESULT_outputs[405]),
        .RESULT_406(RESULT_outputs[406]),
        .RESULT_407(RESULT_outputs[407]),
        .RESULT_408(RESULT_outputs[408]),
        .RESULT_409(RESULT_outputs[409]),
        .RESULT_410(RESULT_outputs[410]),
        .RESULT_411(RESULT_outputs[411]),
        .RESULT_412(RESULT_outputs[412]),
        .RESULT_413(RESULT_outputs[413]),
        .RESULT_414(RESULT_outputs[414]),
        .RESULT_415(RESULT_outputs[415]),
        .RESULT_416(RESULT_outputs[416]),
        .RESULT_417(RESULT_outputs[417]),
        .RESULT_418(RESULT_outputs[418]),
        .RESULT_419(RESULT_outputs[419]),
        .RESULT_420(RESULT_outputs[420]),
        .RESULT_421(RESULT_outputs[421]),
        .RESULT_422(RESULT_outputs[422]),
        .RESULT_423(RESULT_outputs[423]),
        .RESULT_424(RESULT_outputs[424]),
        .RESULT_425(RESULT_outputs[425]),
        .RESULT_426(RESULT_outputs[426]),
        .RESULT_427(RESULT_outputs[427]),
        .RESULT_428(RESULT_outputs[428]),
        .RESULT_429(RESULT_outputs[429]),
        .RESULT_430(RESULT_outputs[430]),
        .RESULT_431(RESULT_outputs[431]),
        .RESULT_432(RESULT_outputs[432]),
        .RESULT_433(RESULT_outputs[433]),
        .RESULT_434(RESULT_outputs[434]),
        .RESULT_435(RESULT_outputs[435]),
        .RESULT_436(RESULT_outputs[436]),
        .RESULT_437(RESULT_outputs[437]),
        .RESULT_438(RESULT_outputs[438]),
        .RESULT_439(RESULT_outputs[439]),
        .RESULT_440(RESULT_outputs[440]),
        .RESULT_441(RESULT_outputs[441]),
        .RESULT_442(RESULT_outputs[442]),
        .RESULT_443(RESULT_outputs[443]),
        .RESULT_444(RESULT_outputs[444]),
        .RESULT_445(RESULT_outputs[445]),
        .RESULT_446(RESULT_outputs[446]),
        .RESULT_447(RESULT_outputs[447]),
        .RESULT_448(RESULT_outputs[448]),
        .RESULT_449(RESULT_outputs[449]),
        .RESULT_450(RESULT_outputs[450]),
        .RESULT_451(RESULT_outputs[451]),
        .RESULT_452(RESULT_outputs[452]),
        .RESULT_453(RESULT_outputs[453]),
        .RESULT_454(RESULT_outputs[454]),
        .RESULT_455(RESULT_outputs[455]),
        .RESULT_456(RESULT_outputs[456]),
        .RESULT_457(RESULT_outputs[457]),
        .RESULT_458(RESULT_outputs[458]),
        .RESULT_459(RESULT_outputs[459]),
        .RESULT_460(RESULT_outputs[460]),
        .RESULT_461(RESULT_outputs[461]),
        .RESULT_462(RESULT_outputs[462]),
        .RESULT_463(RESULT_outputs[463]),
        .RESULT_464(RESULT_outputs[464]),
        .RESULT_465(RESULT_outputs[465]),
        .RESULT_466(RESULT_outputs[466]),
        .RESULT_467(RESULT_outputs[467]),
        .RESULT_468(RESULT_outputs[468]),
        .RESULT_469(RESULT_outputs[469]),
        .RESULT_470(RESULT_outputs[470]),
        .RESULT_471(RESULT_outputs[471]),
        .RESULT_472(RESULT_outputs[472]),
        .RESULT_473(RESULT_outputs[473]),
        .RESULT_474(RESULT_outputs[474]),
        .RESULT_475(RESULT_outputs[475]),
        .RESULT_476(RESULT_outputs[476]),
        .RESULT_477(RESULT_outputs[477]),
        .RESULT_478(RESULT_outputs[478]),
        .RESULT_479(RESULT_outputs[479]),
        .RESULT_480(RESULT_outputs[480]),
        .RESULT_481(RESULT_outputs[481]),
        .RESULT_482(RESULT_outputs[482]),
        .RESULT_483(RESULT_outputs[483]),
        .RESULT_484(RESULT_outputs[484]),
        .RESULT_485(RESULT_outputs[485]),
        .RESULT_486(RESULT_outputs[486]),
        .RESULT_487(RESULT_outputs[487]),
        .RESULT_488(RESULT_outputs[488]),
        .RESULT_489(RESULT_outputs[489]),
        .RESULT_490(RESULT_outputs[490]),
        .RESULT_491(RESULT_outputs[491]),
        .RESULT_492(RESULT_outputs[492]),
        .RESULT_493(RESULT_outputs[493]),
        .RESULT_494(RESULT_outputs[494]),
        .RESULT_495(RESULT_outputs[495]),
        .RESULT_496(RESULT_outputs[496]),
        .RESULT_497(RESULT_outputs[497]),
        .RESULT_498(RESULT_outputs[498]),
        .RESULT_499(RESULT_outputs[499]),
        .RESULT_500(RESULT_outputs[500]),
        .RESULT_501(RESULT_outputs[501]),
        .RESULT_502(RESULT_outputs[502]),
        .RESULT_503(RESULT_outputs[503]),
        .RESULT_504(RESULT_outputs[504]),
        .RESULT_505(RESULT_outputs[505]),
        .RESULT_506(RESULT_outputs[506]),
        .RESULT_507(RESULT_outputs[507]),
        .RESULT_508(RESULT_outputs[508]),
        .RESULT_509(RESULT_outputs[509]),
        .RESULT_510(RESULT_outputs[510]),
        .RESULT_511(RESULT_outputs[511]),
        .RESULT_512(RESULT_outputs[512]),
        .RESULT_513(RESULT_outputs[513]),
        .RESULT_514(RESULT_outputs[514]),
        .RESULT_515(RESULT_outputs[515]),
        .RESULT_516(RESULT_outputs[516]),
        .RESULT_517(RESULT_outputs[517]),
        .RESULT_518(RESULT_outputs[518]),
        .RESULT_519(RESULT_outputs[519]),
        .RESULT_520(RESULT_outputs[520]),
        .RESULT_521(RESULT_outputs[521]),
        .RESULT_522(RESULT_outputs[522]),
        .RESULT_523(RESULT_outputs[523]),
        .RESULT_524(RESULT_outputs[524]),
        .RESULT_525(RESULT_outputs[525]),
        .RESULT_526(RESULT_outputs[526]),
        .RESULT_527(RESULT_outputs[527]),
        .RESULT_528(RESULT_outputs[528]),
        .RESULT_529(RESULT_outputs[529]),
        .RESULT_530(RESULT_outputs[530]),
        .RESULT_531(RESULT_outputs[531]),
        .RESULT_532(RESULT_outputs[532]),
        .RESULT_533(RESULT_outputs[533]),
        .RESULT_534(RESULT_outputs[534]),
        .RESULT_535(RESULT_outputs[535]),
        .RESULT_536(RESULT_outputs[536]),
        .RESULT_537(RESULT_outputs[537]),
        .RESULT_538(RESULT_outputs[538]),
        .RESULT_539(RESULT_outputs[539]),
        .RESULT_540(RESULT_outputs[540]),
        .RESULT_541(RESULT_outputs[541]),
        .RESULT_542(RESULT_outputs[542]),
        .RESULT_543(RESULT_outputs[543]),
        .RESULT_544(RESULT_outputs[544]),
        .RESULT_545(RESULT_outputs[545]),
        .RESULT_546(RESULT_outputs[546]),
        .RESULT_547(RESULT_outputs[547]),
        .RESULT_548(RESULT_outputs[548]),
        .RESULT_549(RESULT_outputs[549]),
        .RESULT_550(RESULT_outputs[550]),
        .RESULT_551(RESULT_outputs[551]),
        .RESULT_552(RESULT_outputs[552]),
        .RESULT_553(RESULT_outputs[553]),
        .RESULT_554(RESULT_outputs[554]),
        .RESULT_555(RESULT_outputs[555]),
        .RESULT_556(RESULT_outputs[556]),
        .RESULT_557(RESULT_outputs[557]),
        .RESULT_558(RESULT_outputs[558]),
        .RESULT_559(RESULT_outputs[559]),
        .RESULT_560(RESULT_outputs[560]),
        .RESULT_561(RESULT_outputs[561]),
        .RESULT_562(RESULT_outputs[562]),
        .RESULT_563(RESULT_outputs[563]),
        .RESULT_564(RESULT_outputs[564]),
        .RESULT_565(RESULT_outputs[565]),
        .RESULT_566(RESULT_outputs[566]),
        .RESULT_567(RESULT_outputs[567]),
        .RESULT_568(RESULT_outputs[568]),
        .RESULT_569(RESULT_outputs[569]),
        .RESULT_570(RESULT_outputs[570]),
        .RESULT_571(RESULT_outputs[571]),
        .RESULT_572(RESULT_outputs[572]),
        .RESULT_573(RESULT_outputs[573]),
        .RESULT_574(RESULT_outputs[574]),
        .RESULT_575(RESULT_outputs[575]),
        .RESULT_576(RESULT_outputs[576]),
        .RESULT_577(RESULT_outputs[577]),
        .RESULT_578(RESULT_outputs[578]),
        .RESULT_579(RESULT_outputs[579]),
        .RESULT_580(RESULT_outputs[580]),
        .RESULT_581(RESULT_outputs[581]),
        .RESULT_582(RESULT_outputs[582]),
        .RESULT_583(RESULT_outputs[583]),
        .RESULT_584(RESULT_outputs[584]),
        .RESULT_585(RESULT_outputs[585]),
        .RESULT_586(RESULT_outputs[586]),
        .RESULT_587(RESULT_outputs[587]),
        .RESULT_588(RESULT_outputs[588]),
        .RESULT_589(RESULT_outputs[589]),
        .RESULT_590(RESULT_outputs[590]),
        .RESULT_591(RESULT_outputs[591]),
        .RESULT_592(RESULT_outputs[592]),
        .RESULT_593(RESULT_outputs[593]),
        .RESULT_594(RESULT_outputs[594]),
        .RESULT_595(RESULT_outputs[595]),
        .RESULT_596(RESULT_outputs[596]),
        .RESULT_597(RESULT_outputs[597]),
        .RESULT_598(RESULT_outputs[598]),
        .RESULT_599(RESULT_outputs[599]),
        .RESULT_600(RESULT_outputs[600]),
        .RESULT_601(RESULT_outputs[601]),
        .RESULT_602(RESULT_outputs[602]),
        .RESULT_603(RESULT_outputs[603]),
        .RESULT_604(RESULT_outputs[604]),
        .RESULT_605(RESULT_outputs[605]),
        .RESULT_606(RESULT_outputs[606]),
        .RESULT_607(RESULT_outputs[607]),
        .RESULT_608(RESULT_outputs[608]),
        .RESULT_609(RESULT_outputs[609]),
        .RESULT_610(RESULT_outputs[610]),
        .RESULT_611(RESULT_outputs[611]),
        .RESULT_612(RESULT_outputs[612]),
        .RESULT_613(RESULT_outputs[613]),
        .RESULT_614(RESULT_outputs[614]),
        .RESULT_615(RESULT_outputs[615]),
        .RESULT_616(RESULT_outputs[616]),
        .RESULT_617(RESULT_outputs[617]),
        .RESULT_618(RESULT_outputs[618]),
        .RESULT_619(RESULT_outputs[619]),
        .RESULT_620(RESULT_outputs[620]),
        .RESULT_621(RESULT_outputs[621]),
        .RESULT_622(RESULT_outputs[622]),
        .RESULT_623(RESULT_outputs[623]),
        .RESULT_624(RESULT_outputs[624]),
        .RESULT_625(RESULT_outputs[625]),
        .RESULT_626(RESULT_outputs[626]),
        .RESULT_627(RESULT_outputs[627]),
        .RESULT_628(RESULT_outputs[628]),
        .RESULT_629(RESULT_outputs[629]),
        .RESULT_630(RESULT_outputs[630]),
        .RESULT_631(RESULT_outputs[631]),
        .RESULT_632(RESULT_outputs[632]),
        .RESULT_633(RESULT_outputs[633]),
        .RESULT_634(RESULT_outputs[634]),
        .RESULT_635(RESULT_outputs[635]),
        .RESULT_636(RESULT_outputs[636]),
        .RESULT_637(RESULT_outputs[637]),
        .RESULT_638(RESULT_outputs[638]),
        .RESULT_639(RESULT_outputs[639]),
        .RESULT_640(RESULT_outputs[640]),
        .RESULT_641(RESULT_outputs[641]),
        .RESULT_642(RESULT_outputs[642]),
        .RESULT_643(RESULT_outputs[643]),
        .RESULT_644(RESULT_outputs[644]),
        .RESULT_645(RESULT_outputs[645]),
        .RESULT_646(RESULT_outputs[646]),
        .RESULT_647(RESULT_outputs[647]),
        .RESULT_648(RESULT_outputs[648]),
        .RESULT_649(RESULT_outputs[649]),
        .RESULT_650(RESULT_outputs[650]),
        .RESULT_651(RESULT_outputs[651]),
        .RESULT_652(RESULT_outputs[652]),
        .RESULT_653(RESULT_outputs[653]),
        .RESULT_654(RESULT_outputs[654]),
        .RESULT_655(RESULT_outputs[655]),
        .RESULT_656(RESULT_outputs[656]),
        .RESULT_657(RESULT_outputs[657]),
        .RESULT_658(RESULT_outputs[658]),
        .RESULT_659(RESULT_outputs[659]),
        .RESULT_660(RESULT_outputs[660]),
        .RESULT_661(RESULT_outputs[661]),
        .RESULT_662(RESULT_outputs[662]),
        .RESULT_663(RESULT_outputs[663]),
        .RESULT_664(RESULT_outputs[664]),
        .RESULT_665(RESULT_outputs[665]),
        .RESULT_666(RESULT_outputs[666]),
        .RESULT_667(RESULT_outputs[667]),
        .RESULT_668(RESULT_outputs[668]),
        .RESULT_669(RESULT_outputs[669]),
        .RESULT_670(RESULT_outputs[670]),
        .RESULT_671(RESULT_outputs[671]),
        .RESULT_672(RESULT_outputs[672]),
        .RESULT_673(RESULT_outputs[673]),
        .RESULT_674(RESULT_outputs[674]),
        .RESULT_675(RESULT_outputs[675]),
        .RESULT_676(RESULT_outputs[676]),
        .RESULT_677(RESULT_outputs[677]),
        .RESULT_678(RESULT_outputs[678]),
        .RESULT_679(RESULT_outputs[679]),
        .RESULT_680(RESULT_outputs[680]),
        .RESULT_681(RESULT_outputs[681]),
        .RESULT_682(RESULT_outputs[682]),
        .RESULT_683(RESULT_outputs[683]),
        .RESULT_684(RESULT_outputs[684]),
        .RESULT_685(RESULT_outputs[685]),
        .RESULT_686(RESULT_outputs[686]),
        .RESULT_687(RESULT_outputs[687]),
        .RESULT_688(RESULT_outputs[688]),
        .RESULT_689(RESULT_outputs[689]),
        .RESULT_690(RESULT_outputs[690]),
        .RESULT_691(RESULT_outputs[691]),
        .RESULT_692(RESULT_outputs[692]),
        .RESULT_693(RESULT_outputs[693]),
        .RESULT_694(RESULT_outputs[694]),
        .RESULT_695(RESULT_outputs[695]),
        .RESULT_696(RESULT_outputs[696]),
        .RESULT_697(RESULT_outputs[697]),
        .RESULT_698(RESULT_outputs[698]),
        .RESULT_699(RESULT_outputs[699]),
        .RESULT_700(RESULT_outputs[700]),
        .RESULT_701(RESULT_outputs[701]),
        .RESULT_702(RESULT_outputs[702]),
        .RESULT_703(RESULT_outputs[703]),
        .RESULT_704(RESULT_outputs[704]),
        .RESULT_705(RESULT_outputs[705]),
        .RESULT_706(RESULT_outputs[706]),
        .RESULT_707(RESULT_outputs[707]),
        .RESULT_708(RESULT_outputs[708]),
        .RESULT_709(RESULT_outputs[709]),
        .RESULT_710(RESULT_outputs[710]),
        .RESULT_711(RESULT_outputs[711]),
        .RESULT_712(RESULT_outputs[712]),
        .RESULT_713(RESULT_outputs[713]),
        .RESULT_714(RESULT_outputs[714]),
        .RESULT_715(RESULT_outputs[715]),
        .RESULT_716(RESULT_outputs[716]),
        .RESULT_717(RESULT_outputs[717]),
        .RESULT_718(RESULT_outputs[718]),
        .RESULT_719(RESULT_outputs[719]),
        .RESULT_720(RESULT_outputs[720]),
        .RESULT_721(RESULT_outputs[721]),
        .RESULT_722(RESULT_outputs[722]),
        .RESULT_723(RESULT_outputs[723]),
        .RESULT_724(RESULT_outputs[724]),
        .RESULT_725(RESULT_outputs[725]),
        .RESULT_726(RESULT_outputs[726]),
        .RESULT_727(RESULT_outputs[727]),
        .RESULT_728(RESULT_outputs[728]),
        .RESULT_729(RESULT_outputs[729]),
        .RESULT_730(RESULT_outputs[730]),
        .RESULT_731(RESULT_outputs[731]),
        .RESULT_732(RESULT_outputs[732]),
        .RESULT_733(RESULT_outputs[733]),
        .RESULT_734(RESULT_outputs[734]),
        .RESULT_735(RESULT_outputs[735]),
        .RESULT_736(RESULT_outputs[736]),
        .RESULT_737(RESULT_outputs[737]),
        .RESULT_738(RESULT_outputs[738]),
        .RESULT_739(RESULT_outputs[739]),
        .RESULT_740(RESULT_outputs[740]),
        .RESULT_741(RESULT_outputs[741]),
        .RESULT_742(RESULT_outputs[742]),
        .RESULT_743(RESULT_outputs[743]),
        .RESULT_744(RESULT_outputs[744]),
        .RESULT_745(RESULT_outputs[745]),
        .RESULT_746(RESULT_outputs[746]),
        .RESULT_747(RESULT_outputs[747]),
        .RESULT_748(RESULT_outputs[748]),
        .RESULT_749(RESULT_outputs[749]),
        .RESULT_750(RESULT_outputs[750]),
        .RESULT_751(RESULT_outputs[751]),
        .RESULT_752(RESULT_outputs[752]),
        .RESULT_753(RESULT_outputs[753]),
        .RESULT_754(RESULT_outputs[754]),
        .RESULT_755(RESULT_outputs[755]),
        .RESULT_756(RESULT_outputs[756]),
        .RESULT_757(RESULT_outputs[757]),
        .RESULT_758(RESULT_outputs[758]),
        .RESULT_759(RESULT_outputs[759]),
        .RESULT_760(RESULT_outputs[760]),
        .RESULT_761(RESULT_outputs[761]),
        .RESULT_762(RESULT_outputs[762]),
        .RESULT_763(RESULT_outputs[763]),
        .RESULT_764(RESULT_outputs[764]),
        .RESULT_765(RESULT_outputs[765]),
        .RESULT_766(RESULT_outputs[766]),
        .RESULT_767(RESULT_outputs[767]),
        .RESULT_768(RESULT_outputs[768]),
        .RESULT_769(RESULT_outputs[769]),
        .RESULT_770(RESULT_outputs[770]),
        .RESULT_771(RESULT_outputs[771]),
        .RESULT_772(RESULT_outputs[772]),
        .RESULT_773(RESULT_outputs[773]),
        .RESULT_774(RESULT_outputs[774]),
        .RESULT_775(RESULT_outputs[775]),
        .RESULT_776(RESULT_outputs[776]),
        .RESULT_777(RESULT_outputs[777]),
        .RESULT_778(RESULT_outputs[778]),
        .RESULT_779(RESULT_outputs[779]),
        .RESULT_780(RESULT_outputs[780]),
        .RESULT_781(RESULT_outputs[781]),
        .RESULT_782(RESULT_outputs[782]),
        .RESULT_783(RESULT_outputs[783]),
        .RESULT_784(RESULT_outputs[784]),
        .RESULT_785(RESULT_outputs[785]),
        .RESULT_786(RESULT_outputs[786]),
        .RESULT_787(RESULT_outputs[787]),
        .RESULT_788(RESULT_outputs[788]),
        .RESULT_789(RESULT_outputs[789]),
        .RESULT_790(RESULT_outputs[790]),
        .RESULT_791(RESULT_outputs[791]),
        .RESULT_792(RESULT_outputs[792]),
        .RESULT_793(RESULT_outputs[793]),
        .RESULT_794(RESULT_outputs[794]),
        .RESULT_795(RESULT_outputs[795]),
        .RESULT_796(RESULT_outputs[796]),
        .RESULT_797(RESULT_outputs[797]),
        .RESULT_798(RESULT_outputs[798]),
        .RESULT_799(RESULT_outputs[799]),
        .RESULT_800(RESULT_outputs[800]),
        .RESULT_801(RESULT_outputs[801]),
        .RESULT_802(RESULT_outputs[802]),
        .RESULT_803(RESULT_outputs[803]),
        .RESULT_804(RESULT_outputs[804]),
        .RESULT_805(RESULT_outputs[805]),
        .RESULT_806(RESULT_outputs[806]),
        .RESULT_807(RESULT_outputs[807]),
        .RESULT_808(RESULT_outputs[808]),
        .RESULT_809(RESULT_outputs[809]),
        .RESULT_810(RESULT_outputs[810]),
        .RESULT_811(RESULT_outputs[811]),
        .RESULT_812(RESULT_outputs[812]),
        .RESULT_813(RESULT_outputs[813]),
        .RESULT_814(RESULT_outputs[814]),
        .RESULT_815(RESULT_outputs[815]),
        .RESULT_816(RESULT_outputs[816]),
        .RESULT_817(RESULT_outputs[817]),
        .RESULT_818(RESULT_outputs[818]),
        .RESULT_819(RESULT_outputs[819]),
        .RESULT_820(RESULT_outputs[820]),
        .RESULT_821(RESULT_outputs[821]),
        .RESULT_822(RESULT_outputs[822]),
        .RESULT_823(RESULT_outputs[823]),
        .RESULT_824(RESULT_outputs[824]),
        .RESULT_825(RESULT_outputs[825]),
        .RESULT_826(RESULT_outputs[826]),
        .RESULT_827(RESULT_outputs[827]),
        .RESULT_828(RESULT_outputs[828]),
        .RESULT_829(RESULT_outputs[829]),
        .RESULT_830(RESULT_outputs[830]),
        .RESULT_831(RESULT_outputs[831]),
        .RESULT_832(RESULT_outputs[832]),
        .RESULT_833(RESULT_outputs[833]),
        .RESULT_834(RESULT_outputs[834]),
        .RESULT_835(RESULT_outputs[835]),
        .RESULT_836(RESULT_outputs[836]),
        .RESULT_837(RESULT_outputs[837]),
        .RESULT_838(RESULT_outputs[838]),
        .RESULT_839(RESULT_outputs[839]),
        .RESULT_840(RESULT_outputs[840]),
        .RESULT_841(RESULT_outputs[841]),
        .RESULT_842(RESULT_outputs[842]),
        .RESULT_843(RESULT_outputs[843]),
        .RESULT_844(RESULT_outputs[844]),
        .RESULT_845(RESULT_outputs[845]),
        .RESULT_846(RESULT_outputs[846]),
        .RESULT_847(RESULT_outputs[847]),
        .RESULT_848(RESULT_outputs[848]),
        .RESULT_849(RESULT_outputs[849]),
        .RESULT_850(RESULT_outputs[850]),
        .RESULT_851(RESULT_outputs[851]),
        .RESULT_852(RESULT_outputs[852]),
        .RESULT_853(RESULT_outputs[853]),
        .RESULT_854(RESULT_outputs[854]),
        .RESULT_855(RESULT_outputs[855]),
        .RESULT_856(RESULT_outputs[856]),
        .RESULT_857(RESULT_outputs[857]),
        .RESULT_858(RESULT_outputs[858]),
        .RESULT_859(RESULT_outputs[859]),
        .RESULT_860(RESULT_outputs[860]),
        .RESULT_861(RESULT_outputs[861]),
        .RESULT_862(RESULT_outputs[862]),
        .RESULT_863(RESULT_outputs[863]),
        .RESULT_864(RESULT_outputs[864]),
        .RESULT_865(RESULT_outputs[865]),
        .RESULT_866(RESULT_outputs[866]),
        .RESULT_867(RESULT_outputs[867]),
        .RESULT_868(RESULT_outputs[868]),
        .RESULT_869(RESULT_outputs[869]),
        .RESULT_870(RESULT_outputs[870]),
        .RESULT_871(RESULT_outputs[871]),
        .RESULT_872(RESULT_outputs[872]),
        .RESULT_873(RESULT_outputs[873]),
        .RESULT_874(RESULT_outputs[874]),
        .RESULT_875(RESULT_outputs[875]),
        .RESULT_876(RESULT_outputs[876]),
        .RESULT_877(RESULT_outputs[877]),
        .RESULT_878(RESULT_outputs[878]),
        .RESULT_879(RESULT_outputs[879]),
        .RESULT_880(RESULT_outputs[880]),
        .RESULT_881(RESULT_outputs[881]),
        .RESULT_882(RESULT_outputs[882]),
        .RESULT_883(RESULT_outputs[883]),
        .RESULT_884(RESULT_outputs[884]),
        .RESULT_885(RESULT_outputs[885]),
        .RESULT_886(RESULT_outputs[886]),
        .RESULT_887(RESULT_outputs[887]),
        .RESULT_888(RESULT_outputs[888]),
        .RESULT_889(RESULT_outputs[889]),
        .RESULT_890(RESULT_outputs[890]),
        .RESULT_891(RESULT_outputs[891]),
        .RESULT_892(RESULT_outputs[892]),
        .RESULT_893(RESULT_outputs[893]),
        .RESULT_894(RESULT_outputs[894]),
        .RESULT_895(RESULT_outputs[895])
    );
    initial begin
             $sdf_annotate("./../../../syn/LAB3/outputs/TOP_gate.sdf",dut);
   
   end

    function real fixed_to_real;
        input [15:0] fixed_val;
        input integer decimal_pos;
        begin
            fixed_to_real = $itor($signed(fixed_val)) / (2.0 ** decimal_pos);
        end
    endfunction

    function real calculate_mxint_snr;
        input logic [15:0] fp16_inputs[];
        input logic [15:0] mxint_outputs[];
        integer i;
        real signal_power, noise_power, diff;
        begin
            signal_power = 0.0;
            noise_power = 0.0;
            for (i = 0; i < NUM_INPUTS; i = i + 1) begin
                diff = fixed_to_real(mxint_outputs[i], DECIMAL_N0) - fp16_to_real(fp16_inputs[i]);
                signal_power += fp16_to_real(fp16_inputs[i]) * fp16_to_real(fp16_inputs[i]);
                noise_power += diff * diff;
            end
            calculate_mxint_snr = 10.0 * $log10(signal_power / noise_power);
        end
    endfunction


    function [15:0] real_to_fp16;
        input real value;
        integer exp;
        real frac;
        integer tmp_val;
        reg sign_bit;

        begin
            if (value == 0.0) begin
                real_to_fp16 = 16'b0;
            end else begin
                if (value < 0.0) begin
                    sign_bit = 1;
                    value = -value;
                end else begin
                    sign_bit = 0;
                end

                exp = $floor($ln(value) / $ln(2.0));
                if (exp != -15) begin
                    frac = value / (2.0 ** exp);
                end else begin
                    frac = value / (2.0 ** -14);
                end
                exp = exp + 15;

                if (exp > 31) begin
                    real_to_fp16 = {sign_bit, 5'b11111, 10'b0};
                end else begin
                    if (exp != 0) begin
                        tmp_val = $rtoi((frac - 1.0) * 1024.0);
                    end else begin
                        tmp_val = $rtoi(frac * 1024.0);
                    end
                    real_to_fp16 = {sign_bit, exp[4:0], tmp_val[9:0]};
                end
            end
        end
    endfunction


    function real fp16_to_real;
        input [15:0] fp16_val;
        integer exp;
        real frac;
        begin
            if (fp16_val[14:10] == 5'b11111) begin
                fp16_to_real = (fp16_val[9:0] == 10'b0) ? $bitstoreal({fp16_val[15], 63'b1111111_10000000_00000000_00000000_00000000_00000000_00000000_00000000}) : 0.0;
            end 
            
            else begin
                exp = fp16_val[14:10] - 15;
                if (exp != -15) begin
                    frac = (1.0 + (fp16_val[9:0] / 1024.0));
                    fp16_to_real = ((fp16_val[15] == 1) ? -1.0 : 1.0) * frac * (2.0 ** exp);
                end
                else begin
                    frac = (fp16_val[9:0] / 1024.0);
                    fp16_to_real = ((fp16_val[15] == 1) ? -1.0 : 1.0) * frac * (2.0 ** -14);
                end
            end
        end
    endfunction

    
    function [15:0] fp16_add;
        input [15:0] a, b;
        real a_real, b_real, result_real;
        begin
            a_real = fp16_to_real(a); 
            b_real = fp16_to_real(b);
            result_real = a_real + b_real; 
            fp16_add = real_to_fp16(result_real); 
        end
    endfunction

    
    function [15:0] fp16_sub;
        input [15:0] a, b;
        real a_real, b_real, result_real;
        begin
            a_real = fp16_to_real(a);
            b_real = fp16_to_real(b);
            result_real = a_real - b_real;
            fp16_sub = real_to_fp16(result_real);
        end
    endfunction

    
    function [15:0] fp16_mul;
        input [15:0] a, b;
        real a_real, b_real, result_real;
        begin
            a_real = fp16_to_real(a);
            b_real = fp16_to_real(b); 
            result_real = a_real * b_real; 
            fp16_mul = real_to_fp16(result_real); 
        end
    endfunction


    task generate_inputs;
        integer i;
        begin
            for (i = 0; i < NUM_INPUTS; i = i + 1) begin
                real random_val;
                if ($urandom_range(1, 100) <= 95) begin
                    random_val = ($urandom() % 100000) / 10000.0 - 5.0;
                end else begin
                    if ($urandom_range(0, 1)) begin
                        random_val = ($urandom() % 150000) / 10000.0 - 20.0;
                    end else begin
                        random_val = ($urandom() % 150000) / 10000.0 + 5.0; 
                    end
                end
                inputs[i] = real_to_fp16(random_val); 
            end
        end
    endtask


    task generate_expected;
        input [1:0] operation;
        integer i, j, k, group_size, num_groups, idx1, idx2, output_idx;
        begin
            group_size = 32;
            num_groups = NUM_INPUTS / group_size;
            output_idx = 0; 

            for (i = 0; i < num_groups - 1; i = i + 1) begin
                for (j = i + 1; j < num_groups; j = j + 1) begin 
                    for (k = 0; k < group_size; k = k + 1) begin 
                        idx1 = k + i * group_size; 
                        idx2 = k + j * group_size; 

                        case (operation)
                            2'b00: FP16_expected[output_idx] = fp16_mul(inputs[idx1], inputs[idx2]);
                            2'b01: FP16_expected[output_idx] = fp16_add(inputs[idx1], inputs[idx2]);
                            2'b10: FP16_expected[output_idx] = fp16_sub(inputs[idx1], inputs[idx2]);
                            default: FP16_expected[output_idx] = 16'b0;
                        endcase

                        output_idx = output_idx + 1;
                    end
                end
            end
        end
    endtask


    function real calculate_result_snr;
        input logic [15:0] fp16_expected[];
        input logic [15:0] result_outputs[];
        integer i;
        real signal_power, noise_power, diff, diff1, diff2;
        begin
            signal_power = 0.0;
            noise_power = 0.0;
            for (i = 0; i < NUM_OUTPUTS; i = i + 1) begin
                diff1 = fixed_to_real(result_outputs[i], DECIMAL_N1);
                diff2 = fp16_to_real(fp16_expected[i]);
                diff = diff1 - diff2;
                $display("Iteration: %0d: diff1 = %0f, diff2 = %0f, diff = %0f", i, diff1, diff2, diff);
                signal_power += fp16_to_real(fp16_expected[i]) * fp16_to_real(fp16_expected[i]);
                noise_power += diff * diff;
            end
            calculate_result_snr = 10.0 * $log10(signal_power / noise_power);
        end
    endfunction

    always #10 CLK = ~CLK;

    initial begin

        CLK = 0;
        RSTN = 0;

        log_file = $fopen("simulation_log.txt", "w");
        if (log_file == 0) begin
            $display("Error: Could not open log file.");
            $stop;
        end

        #5 RSTN = 1;
        generate_inputs();

        @(posedge CLK);
        cycle_count_mxint = 0;
        while (!MXINT_outputs[NUM_INPUTS-1]) begin
            @(posedge CLK);
            cycle_count_mxint = cycle_count_mxint + 1;
        end
        mxint_snr = calculate_mxint_snr(inputs, MXINT_outputs);
        $fwrite(log_file, "SNR (MXINT): %0.2f dB\n", mxint_snr);
        $fwrite(log_file, "Clock Cycles (MXINT): %0d\n", cycle_count_mxint);


        calc = 2'b00;
        generate_expected(calc);
        @(posedge CLK);
        cycle_count_mult = 0;
        while (!RESULT_outputs[NUM_OUTPUTS-1]) begin
            @(posedge CLK);
            cycle_count_mult = cycle_count_mult + 1;
        end
        snr_mult = calculate_result_snr(FP16_expected, RESULT_outputs);
        $fwrite(log_file, "SNR (Multiplication): %0.2f dB\n", snr_mult);
        $fwrite(log_file, "Clock Cycles (Multiplication): %0d\n", cycle_count_mult);

        calc = 2'b01;
        generate_expected(calc);
        @(posedge CLK);
        cycle_count_add = 0;
        while (!RESULT_outputs[NUM_OUTPUTS-1]) begin
            @(posedge CLK);
            cycle_count_add = cycle_count_add + 1;
        end
        snr_add = calculate_result_snr(FP16_expected, RESULT_outputs);
        $fwrite(log_file, "SNR (Addition): %0.2f dB\n", snr_add);
        $fwrite(log_file, "Clock Cycles (Addition): %0d\n", cycle_count_add);

        calc = 2'b10;
        generate_expected(calc);
        @(posedge CLK);
        cycle_count_sub = 0;
        while (!RESULT_outputs[NUM_OUTPUTS-1]) begin
            @(posedge CLK);
            cycle_count_sub = cycle_count_sub + 1;
        end
        snr_sub = calculate_result_snr(FP16_expected, RESULT_outputs);
        $fwrite(log_file, "SNR (Subtraction): %0.2f dB\n", snr_sub);
        $fwrite(log_file, "Clock Cycles (Subtraction): %0d\n", cycle_count_sub);

        $fclose(log_file);
        #100
        $finish;
        //$stop;
    end
endmodule