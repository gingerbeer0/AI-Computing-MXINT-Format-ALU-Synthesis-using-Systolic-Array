module TOP
(input CLK,
input RSTN,
input [1:0] calc,
input [15:0] INPUT_0,
input [15:0] INPUT_1,
input [15:0] INPUT_2,
input [15:0] INPUT_3,
input [15:0] INPUT_4,
input [15:0] INPUT_5,
input [15:0] INPUT_6,
input [15:0] INPUT_7,
input [15:0] INPUT_8,
input [15:0] INPUT_9,
input [15:0] INPUT_10,
input [15:0] INPUT_11,
input [15:0] INPUT_12,
input [15:0] INPUT_13,
input [15:0] INPUT_14,
input [15:0] INPUT_15,
input [15:0] INPUT_16,
input [15:0] INPUT_17,
input [15:0] INPUT_18,
input [15:0] INPUT_19,
input [15:0] INPUT_20,
input [15:0] INPUT_21,
input [15:0] INPUT_22,
input [15:0] INPUT_23,
input [15:0] INPUT_24,
input [15:0] INPUT_25,
input [15:0] INPUT_26,
input [15:0] INPUT_27,
input [15:0] INPUT_28,
input [15:0] INPUT_29,
input [15:0] INPUT_30,
input [15:0] INPUT_31,
input [15:0] INPUT_32,
input [15:0] INPUT_33,
input [15:0] INPUT_34,
input [15:0] INPUT_35,
input [15:0] INPUT_36,
input [15:0] INPUT_37,
input [15:0] INPUT_38,
input [15:0] INPUT_39,
input [15:0] INPUT_40,
input [15:0] INPUT_41,
input [15:0] INPUT_42,
input [15:0] INPUT_43,
input [15:0] INPUT_44,
input [15:0] INPUT_45,
input [15:0] INPUT_46,
input [15:0] INPUT_47,
input [15:0] INPUT_48,
input [15:0] INPUT_49,
input [15:0] INPUT_50,
input [15:0] INPUT_51,
input [15:0] INPUT_52,
input [15:0] INPUT_53,
input [15:0] INPUT_54,
input [15:0] INPUT_55,
input [15:0] INPUT_56,
input [15:0] INPUT_57,
input [15:0] INPUT_58,
input [15:0] INPUT_59,
input [15:0] INPUT_60,
input [15:0] INPUT_61,
input [15:0] INPUT_62,
input [15:0] INPUT_63,
input [15:0] INPUT_64,
input [15:0] INPUT_65,
input [15:0] INPUT_66,
input [15:0] INPUT_67,
input [15:0] INPUT_68,
input [15:0] INPUT_69,
input [15:0] INPUT_70,
input [15:0] INPUT_71,
input [15:0] INPUT_72,
input [15:0] INPUT_73,
input [15:0] INPUT_74,
input [15:0] INPUT_75,
input [15:0] INPUT_76,
input [15:0] INPUT_77,
input [15:0] INPUT_78,
input [15:0] INPUT_79,
input [15:0] INPUT_80,
input [15:0] INPUT_81,
input [15:0] INPUT_82,
input [15:0] INPUT_83,
input [15:0] INPUT_84,
input [15:0] INPUT_85,
input [15:0] INPUT_86,
input [15:0] INPUT_87,
input [15:0] INPUT_88,
input [15:0] INPUT_89,
input [15:0] INPUT_90,
input [15:0] INPUT_91,
input [15:0] INPUT_92,
input [15:0] INPUT_93,
input [15:0] INPUT_94,
input [15:0] INPUT_95,
input [15:0] INPUT_96,
input [15:0] INPUT_97,
input [15:0] INPUT_98,
input [15:0] INPUT_99,
input [15:0] INPUT_100,
input [15:0] INPUT_101,
input [15:0] INPUT_102,
input [15:0] INPUT_103,
input [15:0] INPUT_104,
input [15:0] INPUT_105,
input [15:0] INPUT_106,
input [15:0] INPUT_107,
input [15:0] INPUT_108,
input [15:0] INPUT_109,
input [15:0] INPUT_110,
input [15:0] INPUT_111,
input [15:0] INPUT_112,
input [15:0] INPUT_113,
input [15:0] INPUT_114,
input [15:0] INPUT_115,
input [15:0] INPUT_116,
input [15:0] INPUT_117,
input [15:0] INPUT_118,
input [15:0] INPUT_119,
input [15:0] INPUT_120,
input [15:0] INPUT_121,
input [15:0] INPUT_122,
input [15:0] INPUT_123,
input [15:0] INPUT_124,
input [15:0] INPUT_125,
input [15:0] INPUT_126,
input [15:0] INPUT_127,
input [15:0] INPUT_128,
input [15:0] INPUT_129,
input [15:0] INPUT_130,
input [15:0] INPUT_131,
input [15:0] INPUT_132,
input [15:0] INPUT_133,
input [15:0] INPUT_134,
input [15:0] INPUT_135,
input [15:0] INPUT_136,
input [15:0] INPUT_137,
input [15:0] INPUT_138,
input [15:0] INPUT_139,
input [15:0] INPUT_140,
input [15:0] INPUT_141,
input [15:0] INPUT_142,
input [15:0] INPUT_143,
input [15:0] INPUT_144,
input [15:0] INPUT_145,
input [15:0] INPUT_146,
input [15:0] INPUT_147,
input [15:0] INPUT_148,
input [15:0] INPUT_149,
input [15:0] INPUT_150,
input [15:0] INPUT_151,
input [15:0] INPUT_152,
input [15:0] INPUT_153,
input [15:0] INPUT_154,
input [15:0] INPUT_155,
input [15:0] INPUT_156,
input [15:0] INPUT_157,
input [15:0] INPUT_158,
input [15:0] INPUT_159,
input [15:0] INPUT_160,
input [15:0] INPUT_161,
input [15:0] INPUT_162,
input [15:0] INPUT_163,
input [15:0] INPUT_164,
input [15:0] INPUT_165,
input [15:0] INPUT_166,
input [15:0] INPUT_167,
input [15:0] INPUT_168,
input [15:0] INPUT_169,
input [15:0] INPUT_170,
input [15:0] INPUT_171,
input [15:0] INPUT_172,
input [15:0] INPUT_173,
input [15:0] INPUT_174,
input [15:0] INPUT_175,
input [15:0] INPUT_176,
input [15:0] INPUT_177,
input [15:0] INPUT_178,
input [15:0] INPUT_179,
input [15:0] INPUT_180,
input [15:0] INPUT_181,
input [15:0] INPUT_182,
input [15:0] INPUT_183,
input [15:0] INPUT_184,
input [15:0] INPUT_185,
input [15:0] INPUT_186,
input [15:0] INPUT_187,
input [15:0] INPUT_188,
input [15:0] INPUT_189,
input [15:0] INPUT_190,
input [15:0] INPUT_191,
input [15:0] INPUT_192,
input [15:0] INPUT_193,
input [15:0] INPUT_194,
input [15:0] INPUT_195,
input [15:0] INPUT_196,
input [15:0] INPUT_197,
input [15:0] INPUT_198,
input [15:0] INPUT_199,
input [15:0] INPUT_200,
input [15:0] INPUT_201,
input [15:0] INPUT_202,
input [15:0] INPUT_203,
input [15:0] INPUT_204,
input [15:0] INPUT_205,
input [15:0] INPUT_206,
input [15:0] INPUT_207,
input [15:0] INPUT_208,
input [15:0] INPUT_209,
input [15:0] INPUT_210,
input [15:0] INPUT_211,
input [15:0] INPUT_212,
input [15:0] INPUT_213,
input [15:0] INPUT_214,
input [15:0] INPUT_215,
input [15:0] INPUT_216,
input [15:0] INPUT_217,
input [15:0] INPUT_218,
input [15:0] INPUT_219,
input [15:0] INPUT_220,
input [15:0] INPUT_221,
input [15:0] INPUT_222,
input [15:0] INPUT_223,
input [15:0] INPUT_224,
input [15:0] INPUT_225,
input [15:0] INPUT_226,
input [15:0] INPUT_227,
input [15:0] INPUT_228,
input [15:0] INPUT_229,
input [15:0] INPUT_230,
input [15:0] INPUT_231,
input [15:0] INPUT_232,
input [15:0] INPUT_233,
input [15:0] INPUT_234,
input [15:0] INPUT_235,
input [15:0] INPUT_236,
input [15:0] INPUT_237,
input [15:0] INPUT_238,
input [15:0] INPUT_239,
input [15:0] INPUT_240,
input [15:0] INPUT_241,
input [15:0] INPUT_242,
input [15:0] INPUT_243,
input [15:0] INPUT_244,
input [15:0] INPUT_245,
input [15:0] INPUT_246,
input [15:0] INPUT_247,
input [15:0] INPUT_248,
input [15:0] INPUT_249,
input [15:0] INPUT_250,
input [15:0] INPUT_251,
input [15:0] INPUT_252,
input [15:0] INPUT_253,
input [15:0] INPUT_254,
input [15:0] INPUT_255,

output wire [15:0] MXINT_0,
output wire [15:0] MXINT_1,
output wire [15:0] MXINT_2,
output wire [15:0] MXINT_3,
output wire [15:0] MXINT_4,
output wire [15:0] MXINT_5,
output wire [15:0] MXINT_6,
output wire [15:0] MXINT_7,
output wire [15:0] MXINT_8,
output wire [15:0] MXINT_9,
output wire [15:0] MXINT_10,
output wire [15:0] MXINT_11,
output wire [15:0] MXINT_12,
output wire [15:0] MXINT_13,
output wire [15:0] MXINT_14,
output wire [15:0] MXINT_15,
output wire [15:0] MXINT_16,
output wire [15:0] MXINT_17,
output wire [15:0] MXINT_18,
output wire [15:0] MXINT_19,
output wire [15:0] MXINT_20,
output wire [15:0] MXINT_21,
output wire [15:0] MXINT_22,
output wire [15:0] MXINT_23,
output wire [15:0] MXINT_24,
output wire [15:0] MXINT_25,
output wire [15:0] MXINT_26,
output wire [15:0] MXINT_27,
output wire [15:0] MXINT_28,
output wire [15:0] MXINT_29,
output wire [15:0] MXINT_30,
output wire [15:0] MXINT_31,
output wire [15:0] MXINT_32,
output wire [15:0] MXINT_33,
output wire [15:0] MXINT_34,
output wire [15:0] MXINT_35,
output wire [15:0] MXINT_36,
output wire [15:0] MXINT_37,
output wire [15:0] MXINT_38,
output wire [15:0] MXINT_39,
output wire [15:0] MXINT_40,
output wire [15:0] MXINT_41,
output wire [15:0] MXINT_42,
output wire [15:0] MXINT_43,
output wire [15:0] MXINT_44,
output wire [15:0] MXINT_45,
output wire [15:0] MXINT_46,
output wire [15:0] MXINT_47,
output wire [15:0] MXINT_48,
output wire [15:0] MXINT_49,
output wire [15:0] MXINT_50,
output wire [15:0] MXINT_51,
output wire [15:0] MXINT_52,
output wire [15:0] MXINT_53,
output wire [15:0] MXINT_54,
output wire [15:0] MXINT_55,
output wire [15:0] MXINT_56,
output wire [15:0] MXINT_57,
output wire [15:0] MXINT_58,
output wire [15:0] MXINT_59,
output wire [15:0] MXINT_60,
output wire [15:0] MXINT_61,
output wire [15:0] MXINT_62,
output wire [15:0] MXINT_63,
output wire [15:0] MXINT_64,
output wire [15:0] MXINT_65,
output wire [15:0] MXINT_66,
output wire [15:0] MXINT_67,
output wire [15:0] MXINT_68,
output wire [15:0] MXINT_69,
output wire [15:0] MXINT_70,
output wire [15:0] MXINT_71,
output wire [15:0] MXINT_72,
output wire [15:0] MXINT_73,
output wire [15:0] MXINT_74,
output wire [15:0] MXINT_75,
output wire [15:0] MXINT_76,
output wire [15:0] MXINT_77,
output wire [15:0] MXINT_78,
output wire [15:0] MXINT_79,
output wire [15:0] MXINT_80,
output wire [15:0] MXINT_81,
output wire [15:0] MXINT_82,
output wire [15:0] MXINT_83,
output wire [15:0] MXINT_84,
output wire [15:0] MXINT_85,
output wire [15:0] MXINT_86,
output wire [15:0] MXINT_87,
output wire [15:0] MXINT_88,
output wire [15:0] MXINT_89,
output wire [15:0] MXINT_90,
output wire [15:0] MXINT_91,
output wire [15:0] MXINT_92,
output wire [15:0] MXINT_93,
output wire [15:0] MXINT_94,
output wire [15:0] MXINT_95,
output wire [15:0] MXINT_96,
output wire [15:0] MXINT_97,
output wire [15:0] MXINT_98,
output wire [15:0] MXINT_99,
output wire [15:0] MXINT_100,
output wire [15:0] MXINT_101,
output wire [15:0] MXINT_102,
output wire [15:0] MXINT_103,
output wire [15:0] MXINT_104,
output wire [15:0] MXINT_105,
output wire [15:0] MXINT_106,
output wire [15:0] MXINT_107,
output wire [15:0] MXINT_108,
output wire [15:0] MXINT_109,
output wire [15:0] MXINT_110,
output wire [15:0] MXINT_111,
output wire [15:0] MXINT_112,
output wire [15:0] MXINT_113,
output wire [15:0] MXINT_114,
output wire [15:0] MXINT_115,
output wire [15:0] MXINT_116,
output wire [15:0] MXINT_117,
output wire [15:0] MXINT_118,
output wire [15:0] MXINT_119,
output wire [15:0] MXINT_120,
output wire [15:0] MXINT_121,
output wire [15:0] MXINT_122,
output wire [15:0] MXINT_123,
output wire [15:0] MXINT_124,
output wire [15:0] MXINT_125,
output wire [15:0] MXINT_126,
output wire [15:0] MXINT_127,
output wire [15:0] MXINT_128,
output wire [15:0] MXINT_129,
output wire [15:0] MXINT_130,
output wire [15:0] MXINT_131,
output wire [15:0] MXINT_132,
output wire [15:0] MXINT_133,
output wire [15:0] MXINT_134,
output wire [15:0] MXINT_135,
output wire [15:0] MXINT_136,
output wire [15:0] MXINT_137,
output wire [15:0] MXINT_138,
output wire [15:0] MXINT_139,
output wire [15:0] MXINT_140,
output wire [15:0] MXINT_141,
output wire [15:0] MXINT_142,
output wire [15:0] MXINT_143,
output wire [15:0] MXINT_144,
output wire [15:0] MXINT_145,
output wire [15:0] MXINT_146,
output wire [15:0] MXINT_147,
output wire [15:0] MXINT_148,
output wire [15:0] MXINT_149,
output wire [15:0] MXINT_150,
output wire [15:0] MXINT_151,
output wire [15:0] MXINT_152,
output wire [15:0] MXINT_153,
output wire [15:0] MXINT_154,
output wire [15:0] MXINT_155,
output wire [15:0] MXINT_156,
output wire [15:0] MXINT_157,
output wire [15:0] MXINT_158,
output wire [15:0] MXINT_159,
output wire [15:0] MXINT_160,
output wire [15:0] MXINT_161,
output wire [15:0] MXINT_162,
output wire [15:0] MXINT_163,
output wire [15:0] MXINT_164,
output wire [15:0] MXINT_165,
output wire [15:0] MXINT_166,
output wire [15:0] MXINT_167,
output wire [15:0] MXINT_168,
output wire [15:0] MXINT_169,
output wire [15:0] MXINT_170,
output wire [15:0] MXINT_171,
output wire [15:0] MXINT_172,
output wire [15:0] MXINT_173,
output wire [15:0] MXINT_174,
output wire [15:0] MXINT_175,
output wire [15:0] MXINT_176,
output wire [15:0] MXINT_177,
output wire [15:0] MXINT_178,
output wire [15:0] MXINT_179,
output wire [15:0] MXINT_180,
output wire [15:0] MXINT_181,
output wire [15:0] MXINT_182,
output wire [15:0] MXINT_183,
output wire [15:0] MXINT_184,
output wire [15:0] MXINT_185,
output wire [15:0] MXINT_186,
output wire [15:0] MXINT_187,
output wire [15:0] MXINT_188,
output wire [15:0] MXINT_189,
output wire [15:0] MXINT_190,
output wire [15:0] MXINT_191,
output wire [15:0] MXINT_192,
output wire [15:0] MXINT_193,
output wire [15:0] MXINT_194,
output wire [15:0] MXINT_195,
output wire [15:0] MXINT_196,
output wire [15:0] MXINT_197,
output wire [15:0] MXINT_198,
output wire [15:0] MXINT_199,
output wire [15:0] MXINT_200,
output wire [15:0] MXINT_201,
output wire [15:0] MXINT_202,
output wire [15:0] MXINT_203,
output wire [15:0] MXINT_204,
output wire [15:0] MXINT_205,
output wire [15:0] MXINT_206,
output wire [15:0] MXINT_207,
output wire [15:0] MXINT_208,
output wire [15:0] MXINT_209,
output wire [15:0] MXINT_210,
output wire [15:0] MXINT_211,
output wire [15:0] MXINT_212,
output wire [15:0] MXINT_213,
output wire [15:0] MXINT_214,
output wire [15:0] MXINT_215,
output wire [15:0] MXINT_216,
output wire [15:0] MXINT_217,
output wire [15:0] MXINT_218,
output wire [15:0] MXINT_219,
output wire [15:0] MXINT_220,
output wire [15:0] MXINT_221,
output wire [15:0] MXINT_222,
output wire [15:0] MXINT_223,
output wire [15:0] MXINT_224,
output wire [15:0] MXINT_225,
output wire [15:0] MXINT_226,
output wire [15:0] MXINT_227,
output wire [15:0] MXINT_228,
output wire [15:0] MXINT_229,
output wire [15:0] MXINT_230,
output wire [15:0] MXINT_231,
output wire [15:0] MXINT_232,
output wire [15:0] MXINT_233,
output wire [15:0] MXINT_234,
output wire [15:0] MXINT_235,
output wire [15:0] MXINT_236,
output wire [15:0] MXINT_237,
output wire [15:0] MXINT_238,
output wire [15:0] MXINT_239,
output wire [15:0] MXINT_240,
output wire [15:0] MXINT_241,
output wire [15:0] MXINT_242,
output wire [15:0] MXINT_243,
output wire [15:0] MXINT_244,
output wire [15:0] MXINT_245,
output wire [15:0] MXINT_246,
output wire [15:0] MXINT_247,
output wire [15:0] MXINT_248,
output wire [15:0] MXINT_249,
output wire [15:0] MXINT_250,
output wire [15:0] MXINT_251,
output wire [15:0] MXINT_252,
output wire [15:0] MXINT_253,
output wire [15:0] MXINT_254,
output wire [15:0] MXINT_255,

output wire signed [15:0] RESULT_0,
output wire signed [15:0] RESULT_1,
output wire signed [15:0] RESULT_2,
output wire signed [15:0] RESULT_3,
output wire signed [15:0] RESULT_4,
output wire signed [15:0] RESULT_5,
output wire signed [15:0] RESULT_6,
output wire signed [15:0] RESULT_7,
output wire signed [15:0] RESULT_8,
output wire signed [15:0] RESULT_9,
output wire signed [15:0] RESULT_10,
output wire signed [15:0] RESULT_11,
output wire signed [15:0] RESULT_12,
output wire signed [15:0] RESULT_13,
output wire signed [15:0] RESULT_14,
output wire signed [15:0] RESULT_15,
output wire signed [15:0] RESULT_16,
output wire signed [15:0] RESULT_17,
output wire signed [15:0] RESULT_18,
output wire signed [15:0] RESULT_19,
output wire signed [15:0] RESULT_20,
output wire signed [15:0] RESULT_21,
output wire signed [15:0] RESULT_22,
output wire signed [15:0] RESULT_23,
output wire signed [15:0] RESULT_24,
output wire signed [15:0] RESULT_25,
output wire signed [15:0] RESULT_26,
output wire signed [15:0] RESULT_27,
output wire signed [15:0] RESULT_28,
output wire signed [15:0] RESULT_29,
output wire signed [15:0] RESULT_30,
output wire signed [15:0] RESULT_31,
output wire signed [15:0] RESULT_32,
output wire signed [15:0] RESULT_33,
output wire signed [15:0] RESULT_34,
output wire signed [15:0] RESULT_35,
output wire signed [15:0] RESULT_36,
output wire signed [15:0] RESULT_37,
output wire signed [15:0] RESULT_38,
output wire signed [15:0] RESULT_39,
output wire signed [15:0] RESULT_40,
output wire signed [15:0] RESULT_41,
output wire signed [15:0] RESULT_42,
output wire signed [15:0] RESULT_43,
output wire signed [15:0] RESULT_44,
output wire signed [15:0] RESULT_45,
output wire signed [15:0] RESULT_46,
output wire signed [15:0] RESULT_47,
output wire signed [15:0] RESULT_48,
output wire signed [15:0] RESULT_49,
output wire signed [15:0] RESULT_50,
output wire signed [15:0] RESULT_51,
output wire signed [15:0] RESULT_52,
output wire signed [15:0] RESULT_53,
output wire signed [15:0] RESULT_54,
output wire signed [15:0] RESULT_55,
output wire signed [15:0] RESULT_56,
output wire signed [15:0] RESULT_57,
output wire signed [15:0] RESULT_58,
output wire signed [15:0] RESULT_59,
output wire signed [15:0] RESULT_60,
output wire signed [15:0] RESULT_61,
output wire signed [15:0] RESULT_62,
output wire signed [15:0] RESULT_63,
output wire signed [15:0] RESULT_64,
output wire signed [15:0] RESULT_65,
output wire signed [15:0] RESULT_66,
output wire signed [15:0] RESULT_67,
output wire signed [15:0] RESULT_68,
output wire signed [15:0] RESULT_69,
output wire signed [15:0] RESULT_70,
output wire signed [15:0] RESULT_71,
output wire signed [15:0] RESULT_72,
output wire signed [15:0] RESULT_73,
output wire signed [15:0] RESULT_74,
output wire signed [15:0] RESULT_75,
output wire signed [15:0] RESULT_76,
output wire signed [15:0] RESULT_77,
output wire signed [15:0] RESULT_78,
output wire signed [15:0] RESULT_79,
output wire signed [15:0] RESULT_80,
output wire signed [15:0] RESULT_81,
output wire signed [15:0] RESULT_82,
output wire signed [15:0] RESULT_83,
output wire signed [15:0] RESULT_84,
output wire signed [15:0] RESULT_85,
output wire signed [15:0] RESULT_86,
output wire signed [15:0] RESULT_87,
output wire signed [15:0] RESULT_88,
output wire signed [15:0] RESULT_89,
output wire signed [15:0] RESULT_90,
output wire signed [15:0] RESULT_91,
output wire signed [15:0] RESULT_92,
output wire signed [15:0] RESULT_93,
output wire signed [15:0] RESULT_94,
output wire signed [15:0] RESULT_95,
output wire signed [15:0] RESULT_96,
output wire signed [15:0] RESULT_97,
output wire signed [15:0] RESULT_98,
output wire signed [15:0] RESULT_99,
output wire signed [15:0] RESULT_100,
output wire signed [15:0] RESULT_101,
output wire signed [15:0] RESULT_102,
output wire signed [15:0] RESULT_103,
output wire signed [15:0] RESULT_104,
output wire signed [15:0] RESULT_105,
output wire signed [15:0] RESULT_106,
output wire signed [15:0] RESULT_107,
output wire signed [15:0] RESULT_108,
output wire signed [15:0] RESULT_109,
output wire signed [15:0] RESULT_110,
output wire signed [15:0] RESULT_111,
output wire signed [15:0] RESULT_112,
output wire signed [15:0] RESULT_113,
output wire signed [15:0] RESULT_114,
output wire signed [15:0] RESULT_115,
output wire signed [15:0] RESULT_116,
output wire signed [15:0] RESULT_117,
output wire signed [15:0] RESULT_118,
output wire signed [15:0] RESULT_119,
output wire signed [15:0] RESULT_120,
output wire signed [15:0] RESULT_121,
output wire signed [15:0] RESULT_122,
output wire signed [15:0] RESULT_123,
output wire signed [15:0] RESULT_124,
output wire signed [15:0] RESULT_125,
output wire signed [15:0] RESULT_126,
output wire signed [15:0] RESULT_127,
output wire signed [15:0] RESULT_128,
output wire signed [15:0] RESULT_129,
output wire signed [15:0] RESULT_130,
output wire signed [15:0] RESULT_131,
output wire signed [15:0] RESULT_132,
output wire signed [15:0] RESULT_133,
output wire signed [15:0] RESULT_134,
output wire signed [15:0] RESULT_135,
output wire signed [15:0] RESULT_136,
output wire signed [15:0] RESULT_137,
output wire signed [15:0] RESULT_138,
output wire signed [15:0] RESULT_139,
output wire signed [15:0] RESULT_140,
output wire signed [15:0] RESULT_141,
output wire signed [15:0] RESULT_142,
output wire signed [15:0] RESULT_143,
output wire signed [15:0] RESULT_144,
output wire signed [15:0] RESULT_145,
output wire signed [15:0] RESULT_146,
output wire signed [15:0] RESULT_147,
output wire signed [15:0] RESULT_148,
output wire signed [15:0] RESULT_149,
output wire signed [15:0] RESULT_150,
output wire signed [15:0] RESULT_151,
output wire signed [15:0] RESULT_152,
output wire signed [15:0] RESULT_153,
output wire signed [15:0] RESULT_154,
output wire signed [15:0] RESULT_155,
output wire signed [15:0] RESULT_156,
output wire signed [15:0] RESULT_157,
output wire signed [15:0] RESULT_158,
output wire signed [15:0] RESULT_159,
output wire signed [15:0] RESULT_160,
output wire signed [15:0] RESULT_161,
output wire signed [15:0] RESULT_162,
output wire signed [15:0] RESULT_163,
output wire signed [15:0] RESULT_164,
output wire signed [15:0] RESULT_165,
output wire signed [15:0] RESULT_166,
output wire signed [15:0] RESULT_167,
output wire signed [15:0] RESULT_168,
output wire signed [15:0] RESULT_169,
output wire signed [15:0] RESULT_170,
output wire signed [15:0] RESULT_171,
output wire signed [15:0] RESULT_172,
output wire signed [15:0] RESULT_173,
output wire signed [15:0] RESULT_174,
output wire signed [15:0] RESULT_175,
output wire signed [15:0] RESULT_176,
output wire signed [15:0] RESULT_177,
output wire signed [15:0] RESULT_178,
output wire signed [15:0] RESULT_179,
output wire signed [15:0] RESULT_180,
output wire signed [15:0] RESULT_181,
output wire signed [15:0] RESULT_182,
output wire signed [15:0] RESULT_183,
output wire signed [15:0] RESULT_184,
output wire signed [15:0] RESULT_185,
output wire signed [15:0] RESULT_186,
output wire signed [15:0] RESULT_187,
output wire signed [15:0] RESULT_188,
output wire signed [15:0] RESULT_189,
output wire signed [15:0] RESULT_190,
output wire signed [15:0] RESULT_191,
output wire signed [15:0] RESULT_192,
output wire signed [15:0] RESULT_193,
output wire signed [15:0] RESULT_194,
output wire signed [15:0] RESULT_195,
output wire signed [15:0] RESULT_196,
output wire signed [15:0] RESULT_197,
output wire signed [15:0] RESULT_198,
output wire signed [15:0] RESULT_199,
output wire signed [15:0] RESULT_200,
output wire signed [15:0] RESULT_201,
output wire signed [15:0] RESULT_202,
output wire signed [15:0] RESULT_203,
output wire signed [15:0] RESULT_204,
output wire signed [15:0] RESULT_205,
output wire signed [15:0] RESULT_206,
output wire signed [15:0] RESULT_207,
output wire signed [15:0] RESULT_208,
output wire signed [15:0] RESULT_209,
output wire signed [15:0] RESULT_210,
output wire signed [15:0] RESULT_211,
output wire signed [15:0] RESULT_212,
output wire signed [15:0] RESULT_213,
output wire signed [15:0] RESULT_214,
output wire signed [15:0] RESULT_215,
output wire signed [15:0] RESULT_216,
output wire signed [15:0] RESULT_217,
output wire signed [15:0] RESULT_218,
output wire signed [15:0] RESULT_219,
output wire signed [15:0] RESULT_220,
output wire signed [15:0] RESULT_221,
output wire signed [15:0] RESULT_222,
output wire signed [15:0] RESULT_223,
output wire signed [15:0] RESULT_224,
output wire signed [15:0] RESULT_225,
output wire signed [15:0] RESULT_226,
output wire signed [15:0] RESULT_227,
output wire signed [15:0] RESULT_228,
output wire signed [15:0] RESULT_229,
output wire signed [15:0] RESULT_230,
output wire signed [15:0] RESULT_231,
output wire signed [15:0] RESULT_232,
output wire signed [15:0] RESULT_233,
output wire signed [15:0] RESULT_234,
output wire signed [15:0] RESULT_235,
output wire signed [15:0] RESULT_236,
output wire signed [15:0] RESULT_237,
output wire signed [15:0] RESULT_238,
output wire signed [15:0] RESULT_239,
output wire signed [15:0] RESULT_240,
output wire signed [15:0] RESULT_241,
output wire signed [15:0] RESULT_242,
output wire signed [15:0] RESULT_243,
output wire signed [15:0] RESULT_244,
output wire signed [15:0] RESULT_245,
output wire signed [15:0] RESULT_246,
output wire signed [15:0] RESULT_247,
output wire signed [15:0] RESULT_248,
output wire signed [15:0] RESULT_249,
output wire signed [15:0] RESULT_250,
output wire signed [15:0] RESULT_251,
output wire signed [15:0] RESULT_252,
output wire signed [15:0] RESULT_253,
output wire signed [15:0] RESULT_254,
output wire signed [15:0] RESULT_255,
output wire signed [15:0] RESULT_256,
output wire signed [15:0] RESULT_257,
output wire signed [15:0] RESULT_258,
output wire signed [15:0] RESULT_259,
output wire signed [15:0] RESULT_260,
output wire signed [15:0] RESULT_261,
output wire signed [15:0] RESULT_262,
output wire signed [15:0] RESULT_263,
output wire signed [15:0] RESULT_264,
output wire signed [15:0] RESULT_265,
output wire signed [15:0] RESULT_266,
output wire signed [15:0] RESULT_267,
output wire signed [15:0] RESULT_268,
output wire signed [15:0] RESULT_269,
output wire signed [15:0] RESULT_270,
output wire signed [15:0] RESULT_271,
output wire signed [15:0] RESULT_272,
output wire signed [15:0] RESULT_273,
output wire signed [15:0] RESULT_274,
output wire signed [15:0] RESULT_275,
output wire signed [15:0] RESULT_276,
output wire signed [15:0] RESULT_277,
output wire signed [15:0] RESULT_278,
output wire signed [15:0] RESULT_279,
output wire signed [15:0] RESULT_280,
output wire signed [15:0] RESULT_281,
output wire signed [15:0] RESULT_282,
output wire signed [15:0] RESULT_283,
output wire signed [15:0] RESULT_284,
output wire signed [15:0] RESULT_285,
output wire signed [15:0] RESULT_286,
output wire signed [15:0] RESULT_287,
output wire signed [15:0] RESULT_288,
output wire signed [15:0] RESULT_289,
output wire signed [15:0] RESULT_290,
output wire signed [15:0] RESULT_291,
output wire signed [15:0] RESULT_292,
output wire signed [15:0] RESULT_293,
output wire signed [15:0] RESULT_294,
output wire signed [15:0] RESULT_295,
output wire signed [15:0] RESULT_296,
output wire signed [15:0] RESULT_297,
output wire signed [15:0] RESULT_298,
output wire signed [15:0] RESULT_299,
output wire signed [15:0] RESULT_300,
output wire signed [15:0] RESULT_301,
output wire signed [15:0] RESULT_302,
output wire signed [15:0] RESULT_303,
output wire signed [15:0] RESULT_304,
output wire signed [15:0] RESULT_305,
output wire signed [15:0] RESULT_306,
output wire signed [15:0] RESULT_307,
output wire signed [15:0] RESULT_308,
output wire signed [15:0] RESULT_309,
output wire signed [15:0] RESULT_310,
output wire signed [15:0] RESULT_311,
output wire signed [15:0] RESULT_312,
output wire signed [15:0] RESULT_313,
output wire signed [15:0] RESULT_314,
output wire signed [15:0] RESULT_315,
output wire signed [15:0] RESULT_316,
output wire signed [15:0] RESULT_317,
output wire signed [15:0] RESULT_318,
output wire signed [15:0] RESULT_319,
output wire signed [15:0] RESULT_320,
output wire signed [15:0] RESULT_321,
output wire signed [15:0] RESULT_322,
output wire signed [15:0] RESULT_323,
output wire signed [15:0] RESULT_324,
output wire signed [15:0] RESULT_325,
output wire signed [15:0] RESULT_326,
output wire signed [15:0] RESULT_327,
output wire signed [15:0] RESULT_328,
output wire signed [15:0] RESULT_329,
output wire signed [15:0] RESULT_330,
output wire signed [15:0] RESULT_331,
output wire signed [15:0] RESULT_332,
output wire signed [15:0] RESULT_333,
output wire signed [15:0] RESULT_334,
output wire signed [15:0] RESULT_335,
output wire signed [15:0] RESULT_336,
output wire signed [15:0] RESULT_337,
output wire signed [15:0] RESULT_338,
output wire signed [15:0] RESULT_339,
output wire signed [15:0] RESULT_340,
output wire signed [15:0] RESULT_341,
output wire signed [15:0] RESULT_342,
output wire signed [15:0] RESULT_343,
output wire signed [15:0] RESULT_344,
output wire signed [15:0] RESULT_345,
output wire signed [15:0] RESULT_346,
output wire signed [15:0] RESULT_347,
output wire signed [15:0] RESULT_348,
output wire signed [15:0] RESULT_349,
output wire signed [15:0] RESULT_350,
output wire signed [15:0] RESULT_351,
output wire signed [15:0] RESULT_352,
output wire signed [15:0] RESULT_353,
output wire signed [15:0] RESULT_354,
output wire signed [15:0] RESULT_355,
output wire signed [15:0] RESULT_356,
output wire signed [15:0] RESULT_357,
output wire signed [15:0] RESULT_358,
output wire signed [15:0] RESULT_359,
output wire signed [15:0] RESULT_360,
output wire signed [15:0] RESULT_361,
output wire signed [15:0] RESULT_362,
output wire signed [15:0] RESULT_363,
output wire signed [15:0] RESULT_364,
output wire signed [15:0] RESULT_365,
output wire signed [15:0] RESULT_366,
output wire signed [15:0] RESULT_367,
output wire signed [15:0] RESULT_368,
output wire signed [15:0] RESULT_369,
output wire signed [15:0] RESULT_370,
output wire signed [15:0] RESULT_371,
output wire signed [15:0] RESULT_372,
output wire signed [15:0] RESULT_373,
output wire signed [15:0] RESULT_374,
output wire signed [15:0] RESULT_375,
output wire signed [15:0] RESULT_376,
output wire signed [15:0] RESULT_377,
output wire signed [15:0] RESULT_378,
output wire signed [15:0] RESULT_379,
output wire signed [15:0] RESULT_380,
output wire signed [15:0] RESULT_381,
output wire signed [15:0] RESULT_382,
output wire signed [15:0] RESULT_383,
output wire signed [15:0] RESULT_384,
output wire signed [15:0] RESULT_385,
output wire signed [15:0] RESULT_386,
output wire signed [15:0] RESULT_387,
output wire signed [15:0] RESULT_388,
output wire signed [15:0] RESULT_389,
output wire signed [15:0] RESULT_390,
output wire signed [15:0] RESULT_391,
output wire signed [15:0] RESULT_392,
output wire signed [15:0] RESULT_393,
output wire signed [15:0] RESULT_394,
output wire signed [15:0] RESULT_395,
output wire signed [15:0] RESULT_396,
output wire signed [15:0] RESULT_397,
output wire signed [15:0] RESULT_398,
output wire signed [15:0] RESULT_399,
output wire signed [15:0] RESULT_400,
output wire signed [15:0] RESULT_401,
output wire signed [15:0] RESULT_402,
output wire signed [15:0] RESULT_403,
output wire signed [15:0] RESULT_404,
output wire signed [15:0] RESULT_405,
output wire signed [15:0] RESULT_406,
output wire signed [15:0] RESULT_407,
output wire signed [15:0] RESULT_408,
output wire signed [15:0] RESULT_409,
output wire signed [15:0] RESULT_410,
output wire signed [15:0] RESULT_411,
output wire signed [15:0] RESULT_412,
output wire signed [15:0] RESULT_413,
output wire signed [15:0] RESULT_414,
output wire signed [15:0] RESULT_415,
output wire signed [15:0] RESULT_416,
output wire signed [15:0] RESULT_417,
output wire signed [15:0] RESULT_418,
output wire signed [15:0] RESULT_419,
output wire signed [15:0] RESULT_420,
output wire signed [15:0] RESULT_421,
output wire signed [15:0] RESULT_422,
output wire signed [15:0] RESULT_423,
output wire signed [15:0] RESULT_424,
output wire signed [15:0] RESULT_425,
output wire signed [15:0] RESULT_426,
output wire signed [15:0] RESULT_427,
output wire signed [15:0] RESULT_428,
output wire signed [15:0] RESULT_429,
output wire signed [15:0] RESULT_430,
output wire signed [15:0] RESULT_431,
output wire signed [15:0] RESULT_432,
output wire signed [15:0] RESULT_433,
output wire signed [15:0] RESULT_434,
output wire signed [15:0] RESULT_435,
output wire signed [15:0] RESULT_436,
output wire signed [15:0] RESULT_437,
output wire signed [15:0] RESULT_438,
output wire signed [15:0] RESULT_439,
output wire signed [15:0] RESULT_440,
output wire signed [15:0] RESULT_441,
output wire signed [15:0] RESULT_442,
output wire signed [15:0] RESULT_443,
output wire signed [15:0] RESULT_444,
output wire signed [15:0] RESULT_445,
output wire signed [15:0] RESULT_446,
output wire signed [15:0] RESULT_447,
output wire signed [15:0] RESULT_448,
output wire signed [15:0] RESULT_449,
output wire signed [15:0] RESULT_450,
output wire signed [15:0] RESULT_451,
output wire signed [15:0] RESULT_452,
output wire signed [15:0] RESULT_453,
output wire signed [15:0] RESULT_454,
output wire signed [15:0] RESULT_455,
output wire signed [15:0] RESULT_456,
output wire signed [15:0] RESULT_457,
output wire signed [15:0] RESULT_458,
output wire signed [15:0] RESULT_459,
output wire signed [15:0] RESULT_460,
output wire signed [15:0] RESULT_461,
output wire signed [15:0] RESULT_462,
output wire signed [15:0] RESULT_463,
output wire signed [15:0] RESULT_464,
output wire signed [15:0] RESULT_465,
output wire signed [15:0] RESULT_466,
output wire signed [15:0] RESULT_467,
output wire signed [15:0] RESULT_468,
output wire signed [15:0] RESULT_469,
output wire signed [15:0] RESULT_470,
output wire signed [15:0] RESULT_471,
output wire signed [15:0] RESULT_472,
output wire signed [15:0] RESULT_473,
output wire signed [15:0] RESULT_474,
output wire signed [15:0] RESULT_475,
output wire signed [15:0] RESULT_476,
output wire signed [15:0] RESULT_477,
output wire signed [15:0] RESULT_478,
output wire signed [15:0] RESULT_479,
output wire signed [15:0] RESULT_480,
output wire signed [15:0] RESULT_481,
output wire signed [15:0] RESULT_482,
output wire signed [15:0] RESULT_483,
output wire signed [15:0] RESULT_484,
output wire signed [15:0] RESULT_485,
output wire signed [15:0] RESULT_486,
output wire signed [15:0] RESULT_487,
output wire signed [15:0] RESULT_488,
output wire signed [15:0] RESULT_489,
output wire signed [15:0] RESULT_490,
output wire signed [15:0] RESULT_491,
output wire signed [15:0] RESULT_492,
output wire signed [15:0] RESULT_493,
output wire signed [15:0] RESULT_494,
output wire signed [15:0] RESULT_495,
output wire signed [15:0] RESULT_496,
output wire signed [15:0] RESULT_497,
output wire signed [15:0] RESULT_498,
output wire signed [15:0] RESULT_499,
output wire signed [15:0] RESULT_500,
output wire signed [15:0] RESULT_501,
output wire signed [15:0] RESULT_502,
output wire signed [15:0] RESULT_503,
output wire signed [15:0] RESULT_504,
output wire signed [15:0] RESULT_505,
output wire signed [15:0] RESULT_506,
output wire signed [15:0] RESULT_507,
output wire signed [15:0] RESULT_508,
output wire signed [15:0] RESULT_509,
output wire signed [15:0] RESULT_510,
output wire signed [15:0] RESULT_511,
output wire signed [15:0] RESULT_512,
output wire signed [15:0] RESULT_513,
output wire signed [15:0] RESULT_514,
output wire signed [15:0] RESULT_515,
output wire signed [15:0] RESULT_516,
output wire signed [15:0] RESULT_517,
output wire signed [15:0] RESULT_518,
output wire signed [15:0] RESULT_519,
output wire signed [15:0] RESULT_520,
output wire signed [15:0] RESULT_521,
output wire signed [15:0] RESULT_522,
output wire signed [15:0] RESULT_523,
output wire signed [15:0] RESULT_524,
output wire signed [15:0] RESULT_525,
output wire signed [15:0] RESULT_526,
output wire signed [15:0] RESULT_527,
output wire signed [15:0] RESULT_528,
output wire signed [15:0] RESULT_529,
output wire signed [15:0] RESULT_530,
output wire signed [15:0] RESULT_531,
output wire signed [15:0] RESULT_532,
output wire signed [15:0] RESULT_533,
output wire signed [15:0] RESULT_534,
output wire signed [15:0] RESULT_535,
output wire signed [15:0] RESULT_536,
output wire signed [15:0] RESULT_537,
output wire signed [15:0] RESULT_538,
output wire signed [15:0] RESULT_539,
output wire signed [15:0] RESULT_540,
output wire signed [15:0] RESULT_541,
output wire signed [15:0] RESULT_542,
output wire signed [15:0] RESULT_543,
output wire signed [15:0] RESULT_544,
output wire signed [15:0] RESULT_545,
output wire signed [15:0] RESULT_546,
output wire signed [15:0] RESULT_547,
output wire signed [15:0] RESULT_548,
output wire signed [15:0] RESULT_549,
output wire signed [15:0] RESULT_550,
output wire signed [15:0] RESULT_551,
output wire signed [15:0] RESULT_552,
output wire signed [15:0] RESULT_553,
output wire signed [15:0] RESULT_554,
output wire signed [15:0] RESULT_555,
output wire signed [15:0] RESULT_556,
output wire signed [15:0] RESULT_557,
output wire signed [15:0] RESULT_558,
output wire signed [15:0] RESULT_559,
output wire signed [15:0] RESULT_560,
output wire signed [15:0] RESULT_561,
output wire signed [15:0] RESULT_562,
output wire signed [15:0] RESULT_563,
output wire signed [15:0] RESULT_564,
output wire signed [15:0] RESULT_565,
output wire signed [15:0] RESULT_566,
output wire signed [15:0] RESULT_567,
output wire signed [15:0] RESULT_568,
output wire signed [15:0] RESULT_569,
output wire signed [15:0] RESULT_570,
output wire signed [15:0] RESULT_571,
output wire signed [15:0] RESULT_572,
output wire signed [15:0] RESULT_573,
output wire signed [15:0] RESULT_574,
output wire signed [15:0] RESULT_575,
output wire signed [15:0] RESULT_576,
output wire signed [15:0] RESULT_577,
output wire signed [15:0] RESULT_578,
output wire signed [15:0] RESULT_579,
output wire signed [15:0] RESULT_580,
output wire signed [15:0] RESULT_581,
output wire signed [15:0] RESULT_582,
output wire signed [15:0] RESULT_583,
output wire signed [15:0] RESULT_584,
output wire signed [15:0] RESULT_585,
output wire signed [15:0] RESULT_586,
output wire signed [15:0] RESULT_587,
output wire signed [15:0] RESULT_588,
output wire signed [15:0] RESULT_589,
output wire signed [15:0] RESULT_590,
output wire signed [15:0] RESULT_591,
output wire signed [15:0] RESULT_592,
output wire signed [15:0] RESULT_593,
output wire signed [15:0] RESULT_594,
output wire signed [15:0] RESULT_595,
output wire signed [15:0] RESULT_596,
output wire signed [15:0] RESULT_597,
output wire signed [15:0] RESULT_598,
output wire signed [15:0] RESULT_599,
output wire signed [15:0] RESULT_600,
output wire signed [15:0] RESULT_601,
output wire signed [15:0] RESULT_602,
output wire signed [15:0] RESULT_603,
output wire signed [15:0] RESULT_604,
output wire signed [15:0] RESULT_605,
output wire signed [15:0] RESULT_606,
output wire signed [15:0] RESULT_607,
output wire signed [15:0] RESULT_608,
output wire signed [15:0] RESULT_609,
output wire signed [15:0] RESULT_610,
output wire signed [15:0] RESULT_611,
output wire signed [15:0] RESULT_612,
output wire signed [15:0] RESULT_613,
output wire signed [15:0] RESULT_614,
output wire signed [15:0] RESULT_615,
output wire signed [15:0] RESULT_616,
output wire signed [15:0] RESULT_617,
output wire signed [15:0] RESULT_618,
output wire signed [15:0] RESULT_619,
output wire signed [15:0] RESULT_620,
output wire signed [15:0] RESULT_621,
output wire signed [15:0] RESULT_622,
output wire signed [15:0] RESULT_623,
output wire signed [15:0] RESULT_624,
output wire signed [15:0] RESULT_625,
output wire signed [15:0] RESULT_626,
output wire signed [15:0] RESULT_627,
output wire signed [15:0] RESULT_628,
output wire signed [15:0] RESULT_629,
output wire signed [15:0] RESULT_630,
output wire signed [15:0] RESULT_631,
output wire signed [15:0] RESULT_632,
output wire signed [15:0] RESULT_633,
output wire signed [15:0] RESULT_634,
output wire signed [15:0] RESULT_635,
output wire signed [15:0] RESULT_636,
output wire signed [15:0] RESULT_637,
output wire signed [15:0] RESULT_638,
output wire signed [15:0] RESULT_639,
output wire signed [15:0] RESULT_640,
output wire signed [15:0] RESULT_641,
output wire signed [15:0] RESULT_642,
output wire signed [15:0] RESULT_643,
output wire signed [15:0] RESULT_644,
output wire signed [15:0] RESULT_645,
output wire signed [15:0] RESULT_646,
output wire signed [15:0] RESULT_647,
output wire signed [15:0] RESULT_648,
output wire signed [15:0] RESULT_649,
output wire signed [15:0] RESULT_650,
output wire signed [15:0] RESULT_651,
output wire signed [15:0] RESULT_652,
output wire signed [15:0] RESULT_653,
output wire signed [15:0] RESULT_654,
output wire signed [15:0] RESULT_655,
output wire signed [15:0] RESULT_656,
output wire signed [15:0] RESULT_657,
output wire signed [15:0] RESULT_658,
output wire signed [15:0] RESULT_659,
output wire signed [15:0] RESULT_660,
output wire signed [15:0] RESULT_661,
output wire signed [15:0] RESULT_662,
output wire signed [15:0] RESULT_663,
output wire signed [15:0] RESULT_664,
output wire signed [15:0] RESULT_665,
output wire signed [15:0] RESULT_666,
output wire signed [15:0] RESULT_667,
output wire signed [15:0] RESULT_668,
output wire signed [15:0] RESULT_669,
output wire signed [15:0] RESULT_670,
output wire signed [15:0] RESULT_671,
output wire signed [15:0] RESULT_672,
output wire signed [15:0] RESULT_673,
output wire signed [15:0] RESULT_674,
output wire signed [15:0] RESULT_675,
output wire signed [15:0] RESULT_676,
output wire signed [15:0] RESULT_677,
output wire signed [15:0] RESULT_678,
output wire signed [15:0] RESULT_679,
output wire signed [15:0] RESULT_680,
output wire signed [15:0] RESULT_681,
output wire signed [15:0] RESULT_682,
output wire signed [15:0] RESULT_683,
output wire signed [15:0] RESULT_684,
output wire signed [15:0] RESULT_685,
output wire signed [15:0] RESULT_686,
output wire signed [15:0] RESULT_687,
output wire signed [15:0] RESULT_688,
output wire signed [15:0] RESULT_689,
output wire signed [15:0] RESULT_690,
output wire signed [15:0] RESULT_691,
output wire signed [15:0] RESULT_692,
output wire signed [15:0] RESULT_693,
output wire signed [15:0] RESULT_694,
output wire signed [15:0] RESULT_695,
output wire signed [15:0] RESULT_696,
output wire signed [15:0] RESULT_697,
output wire signed [15:0] RESULT_698,
output wire signed [15:0] RESULT_699,
output wire signed [15:0] RESULT_700,
output wire signed [15:0] RESULT_701,
output wire signed [15:0] RESULT_702,
output wire signed [15:0] RESULT_703,
output wire signed [15:0] RESULT_704,
output wire signed [15:0] RESULT_705,
output wire signed [15:0] RESULT_706,
output wire signed [15:0] RESULT_707,
output wire signed [15:0] RESULT_708,
output wire signed [15:0] RESULT_709,
output wire signed [15:0] RESULT_710,
output wire signed [15:0] RESULT_711,
output wire signed [15:0] RESULT_712,
output wire signed [15:0] RESULT_713,
output wire signed [15:0] RESULT_714,
output wire signed [15:0] RESULT_715,
output wire signed [15:0] RESULT_716,
output wire signed [15:0] RESULT_717,
output wire signed [15:0] RESULT_718,
output wire signed [15:0] RESULT_719,
output wire signed [15:0] RESULT_720,
output wire signed [15:0] RESULT_721,
output wire signed [15:0] RESULT_722,
output wire signed [15:0] RESULT_723,
output wire signed [15:0] RESULT_724,
output wire signed [15:0] RESULT_725,
output wire signed [15:0] RESULT_726,
output wire signed [15:0] RESULT_727,
output wire signed [15:0] RESULT_728,
output wire signed [15:0] RESULT_729,
output wire signed [15:0] RESULT_730,
output wire signed [15:0] RESULT_731,
output wire signed [15:0] RESULT_732,
output wire signed [15:0] RESULT_733,
output wire signed [15:0] RESULT_734,
output wire signed [15:0] RESULT_735,
output wire signed [15:0] RESULT_736,
output wire signed [15:0] RESULT_737,
output wire signed [15:0] RESULT_738,
output wire signed [15:0] RESULT_739,
output wire signed [15:0] RESULT_740,
output wire signed [15:0] RESULT_741,
output wire signed [15:0] RESULT_742,
output wire signed [15:0] RESULT_743,
output wire signed [15:0] RESULT_744,
output wire signed [15:0] RESULT_745,
output wire signed [15:0] RESULT_746,
output wire signed [15:0] RESULT_747,
output wire signed [15:0] RESULT_748,
output wire signed [15:0] RESULT_749,
output wire signed [15:0] RESULT_750,
output wire signed [15:0] RESULT_751,
output wire signed [15:0] RESULT_752,
output wire signed [15:0] RESULT_753,
output wire signed [15:0] RESULT_754,
output wire signed [15:0] RESULT_755,
output wire signed [15:0] RESULT_756,
output wire signed [15:0] RESULT_757,
output wire signed [15:0] RESULT_758,
output wire signed [15:0] RESULT_759,
output wire signed [15:0] RESULT_760,
output wire signed [15:0] RESULT_761,
output wire signed [15:0] RESULT_762,
output wire signed [15:0] RESULT_763,
output wire signed [15:0] RESULT_764,
output wire signed [15:0] RESULT_765,
output wire signed [15:0] RESULT_766,
output wire signed [15:0] RESULT_767,
output wire signed [15:0] RESULT_768,
output wire signed [15:0] RESULT_769,
output wire signed [15:0] RESULT_770,
output wire signed [15:0] RESULT_771,
output wire signed [15:0] RESULT_772,
output wire signed [15:0] RESULT_773,
output wire signed [15:0] RESULT_774,
output wire signed [15:0] RESULT_775,
output wire signed [15:0] RESULT_776,
output wire signed [15:0] RESULT_777,
output wire signed [15:0] RESULT_778,
output wire signed [15:0] RESULT_779,
output wire signed [15:0] RESULT_780,
output wire signed [15:0] RESULT_781,
output wire signed [15:0] RESULT_782,
output wire signed [15:0] RESULT_783,
output wire signed [15:0] RESULT_784,
output wire signed [15:0] RESULT_785,
output wire signed [15:0] RESULT_786,
output wire signed [15:0] RESULT_787,
output wire signed [15:0] RESULT_788,
output wire signed [15:0] RESULT_789,
output wire signed [15:0] RESULT_790,
output wire signed [15:0] RESULT_791,
output wire signed [15:0] RESULT_792,
output wire signed [15:0] RESULT_793,
output wire signed [15:0] RESULT_794,
output wire signed [15:0] RESULT_795,
output wire signed [15:0] RESULT_796,
output wire signed [15:0] RESULT_797,
output wire signed [15:0] RESULT_798,
output wire signed [15:0] RESULT_799,
output wire signed [15:0] RESULT_800,
output wire signed [15:0] RESULT_801,
output wire signed [15:0] RESULT_802,
output wire signed [15:0] RESULT_803,
output wire signed [15:0] RESULT_804,
output wire signed [15:0] RESULT_805,
output wire signed [15:0] RESULT_806,
output wire signed [15:0] RESULT_807,
output wire signed [15:0] RESULT_808,
output wire signed [15:0] RESULT_809,
output wire signed [15:0] RESULT_810,
output wire signed [15:0] RESULT_811,
output wire signed [15:0] RESULT_812,
output wire signed [15:0] RESULT_813,
output wire signed [15:0] RESULT_814,
output wire signed [15:0] RESULT_815,
output wire signed [15:0] RESULT_816,
output wire signed [15:0] RESULT_817,
output wire signed [15:0] RESULT_818,
output wire signed [15:0] RESULT_819,
output wire signed [15:0] RESULT_820,
output wire signed [15:0] RESULT_821,
output wire signed [15:0] RESULT_822,
output wire signed [15:0] RESULT_823,
output wire signed [15:0] RESULT_824,
output wire signed [15:0] RESULT_825,
output wire signed [15:0] RESULT_826,
output wire signed [15:0] RESULT_827,
output wire signed [15:0] RESULT_828,
output wire signed [15:0] RESULT_829,
output wire signed [15:0] RESULT_830,
output wire signed [15:0] RESULT_831,
output wire signed [15:0] RESULT_832,
output wire signed [15:0] RESULT_833,
output wire signed [15:0] RESULT_834,
output wire signed [15:0] RESULT_835,
output wire signed [15:0] RESULT_836,
output wire signed [15:0] RESULT_837,
output wire signed [15:0] RESULT_838,
output wire signed [15:0] RESULT_839,
output wire signed [15:0] RESULT_840,
output wire signed [15:0] RESULT_841,
output wire signed [15:0] RESULT_842,
output wire signed [15:0] RESULT_843,
output wire signed [15:0] RESULT_844,
output wire signed [15:0] RESULT_845,
output wire signed [15:0] RESULT_846,
output wire signed [15:0] RESULT_847,
output wire signed [15:0] RESULT_848,
output wire signed [15:0] RESULT_849,
output wire signed [15:0] RESULT_850,
output wire signed [15:0] RESULT_851,
output wire signed [15:0] RESULT_852,
output wire signed [15:0] RESULT_853,
output wire signed [15:0] RESULT_854,
output wire signed [15:0] RESULT_855,
output wire signed [15:0] RESULT_856,
output wire signed [15:0] RESULT_857,
output wire signed [15:0] RESULT_858,
output wire signed [15:0] RESULT_859,
output wire signed [15:0] RESULT_860,
output wire signed [15:0] RESULT_861,
output wire signed [15:0] RESULT_862,
output wire signed [15:0] RESULT_863,
output wire signed [15:0] RESULT_864,
output wire signed [15:0] RESULT_865,
output wire signed [15:0] RESULT_866,
output wire signed [15:0] RESULT_867,
output wire signed [15:0] RESULT_868,
output wire signed [15:0] RESULT_869,
output wire signed [15:0] RESULT_870,
output wire signed [15:0] RESULT_871,
output wire signed [15:0] RESULT_872,
output wire signed [15:0] RESULT_873,
output wire signed [15:0] RESULT_874,
output wire signed [15:0] RESULT_875,
output wire signed [15:0] RESULT_876,
output wire signed [15:0] RESULT_877,
output wire signed [15:0] RESULT_878,
output wire signed [15:0] RESULT_879,
output wire signed [15:0] RESULT_880,
output wire signed [15:0] RESULT_881,
output wire signed [15:0] RESULT_882,
output wire signed [15:0] RESULT_883,
output wire signed [15:0] RESULT_884,
output wire signed [15:0] RESULT_885,
output wire signed [15:0] RESULT_886,
output wire signed [15:0] RESULT_887,
output wire signed [15:0] RESULT_888,
output wire signed [15:0] RESULT_889,
output wire signed [15:0] RESULT_890,
output wire signed [15:0] RESULT_891,
output wire signed [15:0] RESULT_892,
output wire signed [15:0] RESULT_893,
output wire signed [15:0] RESULT_894,
output wire signed [15:0] RESULT_895
);

wire [4:0] shared_exponent0;
wire [4:0] shared_exponent1;
wire [4:0] shared_exponent2;
wire [4:0] shared_exponent3;
wire [4:0] shared_exponent4;
wire [4:0] shared_exponent5;
wire [4:0] shared_exponent6;
wire [4:0] shared_exponent7;

wire [15:0] RESULT_P18;
wire [15:0] RESULT_P17;
wire [15:0] RESULT_P16;
wire [15:0] RESULT_P15;
wire [15:0] RESULT_P14;
wire [15:0] RESULT_P13;
wire [15:0] RESULT_P12;
wire [15:0] RESULT_P28;
wire [15:0] RESULT_P27;
wire [15:0] RESULT_P26;
wire [15:0] RESULT_P25;
wire [15:0] RESULT_P24;
wire [15:0] RESULT_P23;
wire [15:0] RESULT_P38;
wire [15:0] RESULT_P37;
wire [15:0] RESULT_P36;
wire [15:0] RESULT_P35;
wire [15:0] RESULT_P34;
wire [15:0] RESULT_P48;
wire [15:0] RESULT_P47;
wire [15:0] RESULT_P46;
wire [15:0] RESULT_P45;
wire [15:0] RESULT_P58;
wire [15:0] RESULT_P57;
wire [15:0] RESULT_P56;
wire [15:0] RESULT_P68;
wire [15:0] RESULT_P67;
wire [15:0] RESULT_P78;

wire result_enable;
wire alu_enable;

reg enable;
reg alu_enable_reg;

always @(posedge CLK or negedge RSTN) begin
	if (!RSTN) begin
		enable <= 1'b0;
	end else begin
		enable <= 1;
	end
end

always @(posedge CLK or negedge RSTN) begin
	if (!RSTN) begin
		alu_enable_reg <= 1'b0;
	end else begin
		alu_enable_reg <= alu_enable;
	end
end


fp16_to_mxint MX0 (.CLK(CLK), .RSTN(RSTN),.enable(enable), .fp16_in0(INPUT_0), .fp16_in1(INPUT_1), .fp16_in2(INPUT_2), .fp16_in3(INPUT_3), .fp16_in4(INPUT_4), .fp16_in5(INPUT_5), .fp16_in6(INPUT_6), .fp16_in7(INPUT_7), .fp16_in8(INPUT_8), .fp16_in9(INPUT_9), .fp16_in10(INPUT_10), .fp16_in11(INPUT_11), .fp16_in12(INPUT_12), .fp16_in13(INPUT_13), .fp16_in14(INPUT_14), .fp16_in15(INPUT_15), .fp16_in16(INPUT_16),.fp16_in17(INPUT_17), .fp16_in18(INPUT_18), .fp16_in19(INPUT_19), .fp16_in20(INPUT_20), .fp16_in21(INPUT_21), .fp16_in22(INPUT_22),.fp16_in23(INPUT_23),.fp16_in24(INPUT_24),.fp16_in25(INPUT_25),.fp16_in26(INPUT_26),.fp16_in27(INPUT_27),.fp16_in28(INPUT_28),.fp16_in29(INPUT_29),.fp16_in30(INPUT_30),.fp16_in31(INPUT_31), .mxint_res0(MXINT_0),.mxint_res1(MXINT_1),.mxint_res2(MXINT_2),.mxint_res3(MXINT_3),.mxint_res4(MXINT_4),.mxint_res5(MXINT_5),.mxint_res6(MXINT_6),.mxint_res7(MXINT_7),.mxint_res8(MXINT_8),.mxint_res9(MXINT_9),.mxint_res10(MXINT_10),.mxint_res11(MXINT_11),.mxint_res12(MXINT_12),.mxint_res13(MXINT_13),.mxint_res14(MXINT_14),.mxint_res15(MXINT_15),.mxint_res16(MXINT_16),.mxint_res17(MXINT_17),.mxint_res18(MXINT_18),.mxint_res19(MXINT_19),.mxint_res20(MXINT_20),.mxint_res21(MXINT_21),.mxint_res22(MXINT_22),.mxint_res23(MXINT_23),.mxint_res24(MXINT_24),.mxint_res25(MXINT_25),.mxint_res26(MXINT_26),.mxint_res27(MXINT_27),.mxint_res28(MXINT_28),.mxint_res29(MXINT_29),.mxint_res30(MXINT_30), .mxint_res31(MXINT_31), .shared_exponent_out(shared_exponent0));
fp16_to_mxint MX1 (.CLK(CLK), .RSTN(RSTN),.enable(enable), .fp16_in0(INPUT_32), .fp16_in1(INPUT_33), .fp16_in2(INPUT_34), .fp16_in3(INPUT_35), .fp16_in4(INPUT_36), .fp16_in5(INPUT_37), .fp16_in6(INPUT_38), .fp16_in7(INPUT_39), .fp16_in8(INPUT_40), .fp16_in9(INPUT_41), .fp16_in10(INPUT_42), .fp16_in11(INPUT_43), .fp16_in12(INPUT_44), .fp16_in13(INPUT_45), .fp16_in14(INPUT_46), .fp16_in15(INPUT_47), .fp16_in16(INPUT_48),.fp16_in17(INPUT_49), .fp16_in18(INPUT_50), .fp16_in19(INPUT_51), .fp16_in20(INPUT_52), .fp16_in21(INPUT_53), .fp16_in22(INPUT_54),.fp16_in23(INPUT_55),.fp16_in24(INPUT_56),.fp16_in25(INPUT_57),.fp16_in26(INPUT_58),.fp16_in27(INPUT_59),.fp16_in28(INPUT_60),.fp16_in29(INPUT_61),.fp16_in30(INPUT_62),.fp16_in31(INPUT_63), .mxint_res0(MXINT_32),.mxint_res1(MXINT_33),.mxint_res2(MXINT_34),.mxint_res3(MXINT_35),.mxint_res4(MXINT_36),.mxint_res5(MXINT_37),.mxint_res6(MXINT_38),.mxint_res7(MXINT_39),.mxint_res8(MXINT_40),.mxint_res9(MXINT_41),.mxint_res10(MXINT_42),.mxint_res11(MXINT_43),.mxint_res12(MXINT_44),.mxint_res13(MXINT_45),.mxint_res14(MXINT_46),.mxint_res15(MXINT_47),.mxint_res16(MXINT_48),.mxint_res17(MXINT_49),.mxint_res18(MXINT_50),.mxint_res19(MXINT_51),.mxint_res20(MXINT_52),.mxint_res21(MXINT_53),.mxint_res22(MXINT_54),.mxint_res23(MXINT_55),.mxint_res24(MXINT_56),.mxint_res25(MXINT_57),.mxint_res26(MXINT_58),.mxint_res27(MXINT_59),.mxint_res28(MXINT_60),.mxint_res29(MXINT_61),.mxint_res30(MXINT_62), .mxint_res31(MXINT_63), .shared_exponent_out(shared_exponent1));
fp16_to_mxint MX2 (.CLK(CLK), .RSTN(RSTN),.enable(enable), .fp16_in0(INPUT_64), .fp16_in1(INPUT_65), .fp16_in2(INPUT_66), .fp16_in3(INPUT_67), .fp16_in4(INPUT_68), .fp16_in5(INPUT_69), .fp16_in6(INPUT_70), .fp16_in7(INPUT_71), .fp16_in8(INPUT_72), .fp16_in9(INPUT_73), .fp16_in10(INPUT_74), .fp16_in11(INPUT_75), .fp16_in12(INPUT_76), .fp16_in13(INPUT_77), .fp16_in14(INPUT_78), .fp16_in15(INPUT_79), .fp16_in16(INPUT_80),.fp16_in17(INPUT_81), .fp16_in18(INPUT_82), .fp16_in19(INPUT_83), .fp16_in20(INPUT_84), .fp16_in21(INPUT_85), .fp16_in22(INPUT_86),.fp16_in23(INPUT_87),.fp16_in24(INPUT_88),.fp16_in25(INPUT_89),.fp16_in26(INPUT_90),.fp16_in27(INPUT_91),.fp16_in28(INPUT_92),.fp16_in29(INPUT_93),.fp16_in30(INPUT_94),.fp16_in31(INPUT_95), .mxint_res0(MXINT_64),.mxint_res1(MXINT_65),.mxint_res2(MXINT_66),.mxint_res3(MXINT_67),.mxint_res4(MXINT_68),.mxint_res5(MXINT_69),.mxint_res6(MXINT_70),.mxint_res7(MXINT_71),.mxint_res8(MXINT_72),.mxint_res9(MXINT_73),.mxint_res10(MXINT_74),.mxint_res11(MXINT_75),.mxint_res12(MXINT_76),.mxint_res13(MXINT_77),.mxint_res14(MXINT_78),.mxint_res15(MXINT_79),.mxint_res16(MXINT_80),.mxint_res17(MXINT_81),.mxint_res18(MXINT_82),.mxint_res19(MXINT_83),.mxint_res20(MXINT_84),.mxint_res21(MXINT_85),.mxint_res22(MXINT_86),.mxint_res23(MXINT_87),.mxint_res24(MXINT_88),.mxint_res25(MXINT_89),.mxint_res26(MXINT_90),.mxint_res27(MXINT_91),.mxint_res28(MXINT_92),.mxint_res29(MXINT_93),.mxint_res30(MXINT_94), .mxint_res31(MXINT_95), .shared_exponent_out(shared_exponent2));
fp16_to_mxint MX3 (.CLK(CLK), .RSTN(RSTN),.enable(enable), .fp16_in0(INPUT_96), .fp16_in1(INPUT_97), .fp16_in2(INPUT_98), .fp16_in3(INPUT_99), .fp16_in4(INPUT_100), .fp16_in5(INPUT_101), .fp16_in6(INPUT_102), .fp16_in7(INPUT_103), .fp16_in8(INPUT_104), .fp16_in9(INPUT_105), .fp16_in10(INPUT_106), .fp16_in11(INPUT_107), .fp16_in12(INPUT_108), .fp16_in13(INPUT_109), .fp16_in14(INPUT_110), .fp16_in15(INPUT_111), .fp16_in16(INPUT_112),.fp16_in17(INPUT_113), .fp16_in18(INPUT_114), .fp16_in19(INPUT_115), .fp16_in20(INPUT_116), .fp16_in21(INPUT_117), .fp16_in22(INPUT_118),.fp16_in23(INPUT_119),.fp16_in24(INPUT_120),.fp16_in25(INPUT_121),.fp16_in26(INPUT_122),.fp16_in27(INPUT_123),.fp16_in28(INPUT_124),.fp16_in29(INPUT_125),.fp16_in30(INPUT_126),.fp16_in31(INPUT_127), .mxint_res0(MXINT_96),.mxint_res1(MXINT_97),.mxint_res2(MXINT_98),.mxint_res3(MXINT_99),.mxint_res4(MXINT_100),.mxint_res5(MXINT_101),.mxint_res6(MXINT_102),.mxint_res7(MXINT_103),.mxint_res8(MXINT_104),.mxint_res9(MXINT_105),.mxint_res10(MXINT_106),.mxint_res11(MXINT_107),.mxint_res12(MXINT_108),.mxint_res13(MXINT_109),.mxint_res14(MXINT_110),.mxint_res15(MXINT_111),.mxint_res16(MXINT_112),.mxint_res17(MXINT_113),.mxint_res18(MXINT_114),.mxint_res19(MXINT_115),.mxint_res20(MXINT_116),.mxint_res21(MXINT_117),.mxint_res22(MXINT_118),.mxint_res23(MXINT_119),.mxint_res24(MXINT_120),.mxint_res25(MXINT_121),.mxint_res26(MXINT_122),.mxint_res27(MXINT_123),.mxint_res28(MXINT_124),.mxint_res29(MXINT_125),.mxint_res30(MXINT_126),.mxint_res31(MXINT_127), .shared_exponent_out(shared_exponent3));
fp16_to_mxint MX4 (.CLK(CLK), .RSTN(RSTN),.enable(enable), .fp16_in0(INPUT_128), .fp16_in1(INPUT_129), .fp16_in2(INPUT_130), .fp16_in3(INPUT_131), .fp16_in4(INPUT_132), .fp16_in5(INPUT_133), .fp16_in6(INPUT_134), .fp16_in7(INPUT_135), .fp16_in8(INPUT_136), .fp16_in9(INPUT_137), .fp16_in10(INPUT_138), .fp16_in11(INPUT_139), .fp16_in12(INPUT_140), .fp16_in13(INPUT_141), .fp16_in14(INPUT_142), .fp16_in15(INPUT_143), .fp16_in16(INPUT_144),.fp16_in17(INPUT_145), .fp16_in18(INPUT_146), .fp16_in19(INPUT_147), .fp16_in20(INPUT_148), .fp16_in21(INPUT_149), .fp16_in22(INPUT_150),.fp16_in23(INPUT_151),.fp16_in24(INPUT_152),.fp16_in25(INPUT_153),.fp16_in26(INPUT_154),.fp16_in27(INPUT_155),.fp16_in28(INPUT_156),.fp16_in29(INPUT_157),.fp16_in30(INPUT_158),.fp16_in31(INPUT_159), .mxint_res0(MXINT_128),.mxint_res1(MXINT_129),.mxint_res2(MXINT_130),.mxint_res3(MXINT_131),.mxint_res4(MXINT_132),.mxint_res5(MXINT_133),.mxint_res6(MXINT_134),.mxint_res7(MXINT_135),.mxint_res8(MXINT_136),.mxint_res9(MXINT_137),.mxint_res10(MXINT_138),.mxint_res11(MXINT_139),.mxint_res12(MXINT_140),.mxint_res13(MXINT_141),.mxint_res14(MXINT_142),.mxint_res15(MXINT_143),.mxint_res16(MXINT_144),.mxint_res17(MXINT_145),.mxint_res18(MXINT_146),.mxint_res19(MXINT_147),.mxint_res20(MXINT_148),.mxint_res21(MXINT_149),.mxint_res22(MXINT_150),.mxint_res23(MXINT_151),.mxint_res24(MXINT_152),.mxint_res25(MXINT_153),.mxint_res26(MXINT_154),.mxint_res27(MXINT_155),.mxint_res28(MXINT_156),.mxint_res29(MXINT_157),.mxint_res30(MXINT_158), .mxint_res31(MXINT_159), .shared_exponent_out(shared_exponent4));
fp16_to_mxint MX5 (.CLK(CLK), .RSTN(RSTN),.enable(enable), .fp16_in0(INPUT_160), .fp16_in1(INPUT_161), .fp16_in2(INPUT_162), .fp16_in3(INPUT_163), .fp16_in4(INPUT_164), .fp16_in5(INPUT_165), .fp16_in6(INPUT_166), .fp16_in7(INPUT_167), .fp16_in8(INPUT_168), .fp16_in9(INPUT_169), .fp16_in10(INPUT_170), .fp16_in11(INPUT_171), .fp16_in12(INPUT_172), .fp16_in13(INPUT_173), .fp16_in14(INPUT_174), .fp16_in15(INPUT_175), .fp16_in16(INPUT_176),.fp16_in17(INPUT_177), .fp16_in18(INPUT_178), .fp16_in19(INPUT_179), .fp16_in20(INPUT_180), .fp16_in21(INPUT_181), .fp16_in22(INPUT_182),.fp16_in23(INPUT_183),.fp16_in24(INPUT_184),.fp16_in25(INPUT_185),.fp16_in26(INPUT_186),.fp16_in27(INPUT_187),.fp16_in28(INPUT_188),.fp16_in29(INPUT_189),.fp16_in30(INPUT_190),.fp16_in31(INPUT_191), .mxint_res0(MXINT_160),.mxint_res1(MXINT_161),.mxint_res2(MXINT_162),.mxint_res3(MXINT_163),.mxint_res4(MXINT_164),.mxint_res5(MXINT_165),.mxint_res6(MXINT_166),.mxint_res7(MXINT_167),.mxint_res8(MXINT_168),.mxint_res9(MXINT_169),.mxint_res10(MXINT_170),.mxint_res11(MXINT_171),.mxint_res12(MXINT_172),.mxint_res13(MXINT_173),.mxint_res14(MXINT_174),.mxint_res15(MXINT_175),.mxint_res16(MXINT_176),.mxint_res17(MXINT_177),.mxint_res18(MXINT_178),.mxint_res19(MXINT_179),.mxint_res20(MXINT_180),.mxint_res21(MXINT_181),.mxint_res22(MXINT_182),.mxint_res23(MXINT_183),.mxint_res24(MXINT_184),.mxint_res25(MXINT_185),.mxint_res26(MXINT_186),.mxint_res27(MXINT_187),.mxint_res28(MXINT_188),.mxint_res29(MXINT_189),.mxint_res30(MXINT_190), .mxint_res31(MXINT_191), .shared_exponent_out(shared_exponent5));
fp16_to_mxint MX6 (.CLK(CLK), .RSTN(RSTN),.enable(enable), .fp16_in0(INPUT_192), .fp16_in1(INPUT_193), .fp16_in2(INPUT_194), .fp16_in3(INPUT_195), .fp16_in4(INPUT_196), .fp16_in5(INPUT_197), .fp16_in6(INPUT_198), .fp16_in7(INPUT_199), .fp16_in8(INPUT_200), .fp16_in9(INPUT_201), .fp16_in10(INPUT_202), .fp16_in11(INPUT_203), .fp16_in12(INPUT_204), .fp16_in13(INPUT_205), .fp16_in14(INPUT_206), .fp16_in15(INPUT_207), .fp16_in16(INPUT_208),.fp16_in17(INPUT_209), .fp16_in18(INPUT_210), .fp16_in19(INPUT_211), .fp16_in20(INPUT_212), .fp16_in21(INPUT_213), .fp16_in22(INPUT_214),.fp16_in23(INPUT_215),.fp16_in24(INPUT_216),.fp16_in25(INPUT_217),.fp16_in26(INPUT_218),.fp16_in27(INPUT_219),.fp16_in28(INPUT_220),.fp16_in29(INPUT_221),.fp16_in30(INPUT_222),.fp16_in31(INPUT_223), .mxint_res0(MXINT_192),.mxint_res1(MXINT_193),.mxint_res2(MXINT_194),.mxint_res3(MXINT_195),.mxint_res4(MXINT_196),.mxint_res5(MXINT_197),.mxint_res6(MXINT_198),.mxint_res7(MXINT_199),.mxint_res8(MXINT_200),.mxint_res9(MXINT_201),.mxint_res10(MXINT_202),.mxint_res11(MXINT_203),.mxint_res12(MXINT_204),.mxint_res13(MXINT_205),.mxint_res14(MXINT_206),.mxint_res15(MXINT_207),.mxint_res16(MXINT_208),.mxint_res17(MXINT_209),.mxint_res18(MXINT_210),.mxint_res19(MXINT_211),.mxint_res20(MXINT_212),.mxint_res21(MXINT_213),.mxint_res22(MXINT_214),.mxint_res23(MXINT_215),.mxint_res24(MXINT_216),.mxint_res25(MXINT_217),.mxint_res26(MXINT_218),.mxint_res27(MXINT_219),.mxint_res28(MXINT_220),.mxint_res29(MXINT_221),.mxint_res30(MXINT_222), .mxint_res31(MXINT_223), .shared_exponent_out(shared_exponent6));
fp16_to_mxint MX7 (.CLK(CLK), .RSTN(RSTN), .enable(enable),.fp16_in0(INPUT_224), .fp16_in1(INPUT_225), .fp16_in2(INPUT_226), .fp16_in3(INPUT_227), .fp16_in4(INPUT_228), .fp16_in5(INPUT_229), .fp16_in6(INPUT_230), .fp16_in7(INPUT_231), .fp16_in8(INPUT_232), .fp16_in9(INPUT_233), .fp16_in10(INPUT_234), .fp16_in11(INPUT_235), .fp16_in12(INPUT_236), .fp16_in13(INPUT_237), .fp16_in14(INPUT_238), .fp16_in15(INPUT_239), .fp16_in16(INPUT_240),.fp16_in17(INPUT_241), .fp16_in18(INPUT_242), .fp16_in19(INPUT_243), .fp16_in20(INPUT_244), .fp16_in21(INPUT_245), .fp16_in22(INPUT_246),.fp16_in23(INPUT_247),.fp16_in24(INPUT_248),.fp16_in25(INPUT_249),.fp16_in26(INPUT_250),.fp16_in27(INPUT_251),.fp16_in28(INPUT_252),.fp16_in29(INPUT_253),.fp16_in30(INPUT_254),.fp16_in31(INPUT_255), .mxint_res0(MXINT_224),.mxint_res1(MXINT_225),.mxint_res2(MXINT_226),.mxint_res3(MXINT_227),.mxint_res4(MXINT_228),.mxint_res5(MXINT_229),.mxint_res6(MXINT_230),.mxint_res7(MXINT_231),.mxint_res8(MXINT_232),.mxint_res9(MXINT_233),.mxint_res10(MXINT_234),.mxint_res11(MXINT_235),.mxint_res12(MXINT_236),.mxint_res13(MXINT_237),.mxint_res14(MXINT_238),.mxint_res15(MXINT_239),.mxint_res16(MXINT_240),.mxint_res17(MXINT_241),.mxint_res18(MXINT_242),.mxint_res19(MXINT_243),.mxint_res20(MXINT_244),.mxint_res21(MXINT_245),.mxint_res22(MXINT_246),.mxint_res23(MXINT_247),.mxint_res24(MXINT_248),.mxint_res25(MXINT_249),.mxint_res26(MXINT_250),.mxint_res27(MXINT_251),.mxint_res28(MXINT_252),.mxint_res29(MXINT_253),.mxint_res30(MXINT_254), .mxint_res31(MXINT_255), .shared_exponent_out(shared_exponent7), .alu_enable(alu_enable));

stair_array ST1(.CLK(CLK),.RSTN(RSTN),.operation(calc), .enable(alu_enable_reg), .GROUP1_SE(shared_exponent0),.GROUP2_SE(shared_exponent1),.GROUP3_SE(shared_exponent2),.GROUP4_SE(shared_exponent3),.GROUP5_SE(shared_exponent4),.GROUP6_SE(shared_exponent5),.GROUP7_SE(shared_exponent6),.GROUP8_SE(shared_exponent7),.MXINT_0(MXINT_0),.MXINT_1(MXINT_1),.MXINT_2(MXINT_2),.MXINT_3(MXINT_3),.MXINT_4(MXINT_4),.MXINT_5(MXINT_5),.MXINT_6(MXINT_6),.MXINT_7(MXINT_7),.MXINT_8(MXINT_8),.MXINT_9(MXINT_9),.MXINT_10(MXINT_10),.MXINT_11(MXINT_11),.MXINT_12(MXINT_12),.MXINT_13(MXINT_13),.MXINT_14(MXINT_14),.MXINT_15(MXINT_15),.MXINT_16(MXINT_16),.MXINT_17(MXINT_17),.MXINT_18(MXINT_18),.MXINT_19(MXINT_19),.MXINT_20(MXINT_20),.MXINT_21(MXINT_21),.MXINT_22(MXINT_22),.MXINT_23(MXINT_23),.MXINT_24(MXINT_24),.MXINT_25(MXINT_25),.MXINT_26(MXINT_26),.MXINT_27(MXINT_27),.MXINT_28(MXINT_28),.MXINT_29(MXINT_29),.MXINT_30(MXINT_30),.MXINT_31(MXINT_31),.MXINT_32(MXINT_32),.MXINT_33(MXINT_33),.MXINT_34(MXINT_34),.MXINT_35(MXINT_35),.MXINT_36(MXINT_36),.MXINT_37(MXINT_37),.MXINT_38(MXINT_38),.MXINT_39(MXINT_39),.MXINT_40(MXINT_40),.MXINT_41(MXINT_41),.MXINT_42(MXINT_42),.MXINT_43(MXINT_43),.MXINT_44(MXINT_44),.MXINT_45(MXINT_45),.MXINT_46(MXINT_46),.MXINT_47(MXINT_47),.MXINT_48(MXINT_48),.MXINT_49(MXINT_49),.MXINT_50(MXINT_50),.MXINT_51(MXINT_51),.MXINT_52(MXINT_52),.MXINT_53(MXINT_53),.MXINT_54(MXINT_54),.MXINT_55(MXINT_55),.MXINT_56(MXINT_56),.MXINT_57(MXINT_57),.MXINT_58(MXINT_58),.MXINT_59(MXINT_59),.MXINT_60(MXINT_60),.MXINT_61(MXINT_61),.MXINT_62(MXINT_62),.MXINT_63(MXINT_63),.MXINT_64(MXINT_64),.MXINT_65(MXINT_65),.MXINT_66(MXINT_66),.MXINT_67(MXINT_67),.MXINT_68(MXINT_68),.MXINT_69(MXINT_69),.MXINT_70(MXINT_70),.MXINT_71(MXINT_71),.MXINT_72(MXINT_72),.MXINT_73(MXINT_73),.MXINT_74(MXINT_74),.MXINT_75(MXINT_75),.MXINT_76(MXINT_76),.MXINT_77(MXINT_77),.MXINT_78(MXINT_78),.MXINT_79(MXINT_79),.MXINT_80(MXINT_80),.MXINT_81(MXINT_81),.MXINT_82(MXINT_82),.MXINT_83(MXINT_83),.MXINT_84(MXINT_84),.MXINT_85(MXINT_85),.MXINT_86(MXINT_86),.MXINT_87(MXINT_87),.MXINT_88(MXINT_88),.MXINT_89(MXINT_89),.MXINT_90(MXINT_90),.MXINT_91(MXINT_91),.MXINT_92(MXINT_92),.MXINT_93(MXINT_93),.MXINT_94(MXINT_94),.MXINT_95(MXINT_95),.MXINT_96(MXINT_96),.MXINT_97(MXINT_97),.MXINT_98(MXINT_98),.MXINT_99(MXINT_99),.MXINT_100(MXINT_100),.MXINT_101(MXINT_101),.MXINT_102(MXINT_102),.MXINT_103(MXINT_103),.MXINT_104(MXINT_104),.MXINT_105(MXINT_105),.MXINT_106(MXINT_106),.MXINT_107(MXINT_107),.MXINT_108(MXINT_108),.MXINT_109(MXINT_109),.MXINT_110(MXINT_110),.MXINT_111(MXINT_111),.MXINT_112(MXINT_112),.MXINT_113(MXINT_113),.MXINT_114(MXINT_114),.MXINT_115(MXINT_115),.MXINT_116(MXINT_116),.MXINT_117(MXINT_117),.MXINT_118(MXINT_118),.MXINT_119(MXINT_119),.MXINT_120(MXINT_120),.MXINT_121(MXINT_121),.MXINT_122(MXINT_122),.MXINT_123(MXINT_123),.MXINT_124(MXINT_124),.MXINT_125(MXINT_125),.MXINT_126(MXINT_126),.MXINT_127(MXINT_127),.MXINT_128(MXINT_128),.MXINT_129(MXINT_129),.MXINT_130(MXINT_130),.MXINT_131(MXINT_131),.MXINT_132(MXINT_132),.MXINT_133(MXINT_133),.MXINT_134(MXINT_134),.MXINT_135(MXINT_135),.MXINT_136(MXINT_136),.MXINT_137(MXINT_137),.MXINT_138(MXINT_138),.MXINT_139(MXINT_139),.MXINT_140(MXINT_140),.MXINT_141(MXINT_141),.MXINT_142(MXINT_142),.MXINT_143(MXINT_143),.MXINT_144(MXINT_144),.MXINT_145(MXINT_145),.MXINT_146(MXINT_146),.MXINT_147(MXINT_147),.MXINT_148(MXINT_148),.MXINT_149(MXINT_149),.MXINT_150(MXINT_150),.MXINT_151(MXINT_151),.MXINT_152(MXINT_152),.MXINT_153(MXINT_153),.MXINT_154(MXINT_154),.MXINT_155(MXINT_155),.MXINT_156(MXINT_156),.MXINT_157(MXINT_157),.MXINT_158(MXINT_158),.MXINT_159(MXINT_159),.MXINT_160(MXINT_160),.MXINT_161(MXINT_161),.MXINT_162(MXINT_162),.MXINT_163(MXINT_163),.MXINT_164(MXINT_164),.MXINT_165(MXINT_165),.MXINT_166(MXINT_166),.MXINT_167(MXINT_167),.MXINT_168(MXINT_168),.MXINT_169(MXINT_169),.MXINT_170(MXINT_170),.MXINT_171(MXINT_171),.MXINT_172(MXINT_172),.MXINT_173(MXINT_173),.MXINT_174(MXINT_174),.MXINT_175(MXINT_175),.MXINT_176(MXINT_176),.MXINT_177(MXINT_177),.MXINT_178(MXINT_178),.MXINT_179(MXINT_179),.MXINT_180(MXINT_180),.MXINT_181(MXINT_181),.MXINT_182(MXINT_182),.MXINT_183(MXINT_183),.MXINT_184(MXINT_184),.MXINT_185(MXINT_185),.MXINT_186(MXINT_186),.MXINT_187(MXINT_187),.MXINT_188(MXINT_188),.MXINT_189(MXINT_189),.MXINT_190(MXINT_190),.MXINT_191(MXINT_191),.MXINT_192(MXINT_192),.MXINT_193(MXINT_193),.MXINT_194(MXINT_194),.MXINT_195(MXINT_195),.MXINT_196(MXINT_196),.MXINT_197(MXINT_197),.MXINT_198(MXINT_198),.MXINT_199(MXINT_199),.MXINT_200(MXINT_200),.MXINT_201(MXINT_201),.MXINT_202(MXINT_202),.MXINT_203(MXINT_203),.MXINT_204(MXINT_204),.MXINT_205(MXINT_205),.MXINT_206(MXINT_206),.MXINT_207(MXINT_207),.MXINT_208(MXINT_208),.MXINT_209(MXINT_209),.MXINT_210(MXINT_210),.MXINT_211(MXINT_211),.MXINT_212(MXINT_212),.MXINT_213(MXINT_213),.MXINT_214(MXINT_214),.MXINT_215(MXINT_215),.MXINT_216(MXINT_216),.MXINT_217(MXINT_217),.MXINT_218(MXINT_218),.MXINT_219(MXINT_219),.MXINT_220(MXINT_220),.MXINT_221(MXINT_221),.MXINT_222(MXINT_222),.MXINT_223(MXINT_223),.MXINT_224(MXINT_224),.MXINT_225(MXINT_225),.MXINT_226(MXINT_226),.MXINT_227(MXINT_227),.MXINT_228(MXINT_228),.MXINT_229(MXINT_229),.MXINT_230(MXINT_230),.MXINT_231(MXINT_231),.MXINT_232(MXINT_232),.MXINT_233(MXINT_233),.MXINT_234(MXINT_234),.MXINT_235(MXINT_235),.MXINT_236(MXINT_236),.MXINT_237(MXINT_237),.MXINT_238(MXINT_238),.MXINT_239(MXINT_239),.MXINT_240(MXINT_240),.MXINT_241(MXINT_241),.MXINT_242(MXINT_242),.MXINT_243(MXINT_243),.MXINT_244(MXINT_244),.MXINT_245(MXINT_245),.MXINT_246(MXINT_246),.MXINT_247(MXINT_247),.MXINT_248(MXINT_248),.MXINT_249(MXINT_249),.MXINT_250(MXINT_250),.MXINT_251(MXINT_251),.MXINT_252(MXINT_252),.MXINT_253(MXINT_253),.MXINT_254(MXINT_254),.MXINT_255(MXINT_255),.RESULT_P18(RESULT_P18),.RESULT_P17(RESULT_P17),.RESULT_P16(RESULT_P16),.RESULT_P15(RESULT_P15),.RESULT_P14(RESULT_P14),.RESULT_P13(RESULT_P13),.RESULT_P12(RESULT_P12),.RESULT_P28(RESULT_P28),.RESULT_P27(RESULT_P27),.RESULT_P26(RESULT_P26),.RESULT_P25(RESULT_P25),.RESULT_P24(RESULT_P24),.RESULT_P23(RESULT_P23),.RESULT_P38(RESULT_P38),.RESULT_P37(RESULT_P37),.RESULT_P36(RESULT_P36),.RESULT_P35(RESULT_P35),.RESULT_P34(RESULT_P34),.RESULT_P48(RESULT_P48),.RESULT_P47(RESULT_P47),.RESULT_P46(RESULT_P46),.RESULT_P45(RESULT_P45),.RESULT_P58(RESULT_P58),.RESULT_P57(RESULT_P57),.RESULT_P56(RESULT_P56),.RESULT_P68(RESULT_P68),.RESULT_P67(RESULT_P67),.RESULT_P78(RESULT_P78),.result_enable(result_enable));


output_buffer OB (
	.CLK(CLK), .RSTN(RSTN), .result_enable(result_enable),
	.RESULT_P18(RESULT_P18), .RESULT_P17(RESULT_P17), .RESULT_P16(RESULT_P16), .RESULT_P15(RESULT_P15), .RESULT_P14(RESULT_P14), .RESULT_P13(RESULT_P13), .RESULT_P12(RESULT_P12),
	.RESULT_P28(RESULT_P28), .RESULT_P27(RESULT_P27), .RESULT_P26(RESULT_P26), .RESULT_P25(RESULT_P25), .RESULT_P24(RESULT_P24), .RESULT_P23(RESULT_P23),
	.RESULT_P38(RESULT_P38), .RESULT_P37(RESULT_P37), .RESULT_P36(RESULT_P36), .RESULT_P35(RESULT_P35), .RESULT_P34(RESULT_P34),
	.RESULT_P48(RESULT_P48), .RESULT_P47(RESULT_P47), .RESULT_P46(RESULT_P46), .RESULT_P45(RESULT_P45),
	.RESULT_P58(RESULT_P58), .RESULT_P57(RESULT_P57), .RESULT_P56(RESULT_P56),
	.RESULT_P68(RESULT_P68), .RESULT_P67(RESULT_P67), .RESULT_P78(RESULT_P78),
	.RESULT_0(RESULT_0), .RESULT_1(RESULT_1), .RESULT_2(RESULT_2), .RESULT_3(RESULT_3), .RESULT_4(RESULT_4), .RESULT_5(RESULT_5), .RESULT_6(RESULT_6), .RESULT_7(RESULT_7),
	.RESULT_8(RESULT_8), .RESULT_9(RESULT_9), .RESULT_10(RESULT_10), .RESULT_11(RESULT_11), .RESULT_12(RESULT_12), .RESULT_13(RESULT_13), .RESULT_14(RESULT_14), .RESULT_15(RESULT_15),
	.RESULT_16(RESULT_16), .RESULT_17(RESULT_17), .RESULT_18(RESULT_18), .RESULT_19(RESULT_19), .RESULT_20(RESULT_20), .RESULT_21(RESULT_21), .RESULT_22(RESULT_22), .RESULT_23(RESULT_23),
	.RESULT_24(RESULT_24), .RESULT_25(RESULT_25), .RESULT_26(RESULT_26), .RESULT_27(RESULT_27), .RESULT_28(RESULT_28), .RESULT_29(RESULT_29), .RESULT_30(RESULT_30), .RESULT_31(RESULT_31),
	.RESULT_32(RESULT_32), .RESULT_33(RESULT_33), .RESULT_34(RESULT_34), .RESULT_35(RESULT_35), .RESULT_36(RESULT_36), .RESULT_37(RESULT_37), .RESULT_38(RESULT_38), .RESULT_39(RESULT_39),
	.RESULT_40(RESULT_40), .RESULT_41(RESULT_41), .RESULT_42(RESULT_42), .RESULT_43(RESULT_43), .RESULT_44(RESULT_44), .RESULT_45(RESULT_45), .RESULT_46(RESULT_46), .RESULT_47(RESULT_47),
	.RESULT_48(RESULT_48), .RESULT_49(RESULT_49), .RESULT_50(RESULT_50), .RESULT_51(RESULT_51), .RESULT_52(RESULT_52), .RESULT_53(RESULT_53), .RESULT_54(RESULT_54), .RESULT_55(RESULT_55),
	.RESULT_56(RESULT_56), .RESULT_57(RESULT_57), .RESULT_58(RESULT_58), .RESULT_59(RESULT_59), .RESULT_60(RESULT_60), .RESULT_61(RESULT_61), .RESULT_62(RESULT_62), .RESULT_63(RESULT_63),
	.RESULT_64(RESULT_64), .RESULT_65(RESULT_65), .RESULT_66(RESULT_66), .RESULT_67(RESULT_67), .RESULT_68(RESULT_68), .RESULT_69(RESULT_69), .RESULT_70(RESULT_70), .RESULT_71(RESULT_71),
	.RESULT_72(RESULT_72), .RESULT_73(RESULT_73), .RESULT_74(RESULT_74), .RESULT_75(RESULT_75), .RESULT_76(RESULT_76), .RESULT_77(RESULT_77), .RESULT_78(RESULT_78), .RESULT_79(RESULT_79),
	.RESULT_80(RESULT_80), .RESULT_81(RESULT_81), .RESULT_82(RESULT_82), .RESULT_83(RESULT_83), .RESULT_84(RESULT_84), .RESULT_85(RESULT_85), .RESULT_86(RESULT_86), .RESULT_87(RESULT_87),
	.RESULT_88(RESULT_88), .RESULT_89(RESULT_89), .RESULT_90(RESULT_90), .RESULT_91(RESULT_91), .RESULT_92(RESULT_92), .RESULT_93(RESULT_93), .RESULT_94(RESULT_94), .RESULT_95(RESULT_95),
	.RESULT_96(RESULT_96), .RESULT_97(RESULT_97), .RESULT_98(RESULT_98), .RESULT_99(RESULT_99), .RESULT_100(RESULT_100), .RESULT_101(RESULT_101), .RESULT_102(RESULT_102), .RESULT_103(RESULT_103),
	.RESULT_104(RESULT_104), .RESULT_105(RESULT_105), .RESULT_106(RESULT_106), .RESULT_107(RESULT_107), .RESULT_108(RESULT_108), .RESULT_109(RESULT_109), .RESULT_110(RESULT_110), .RESULT_111(RESULT_111),
	.RESULT_112(RESULT_112), .RESULT_113(RESULT_113), .RESULT_114(RESULT_114), .RESULT_115(RESULT_115), .RESULT_116(RESULT_116), .RESULT_117(RESULT_117), .RESULT_118(RESULT_118), .RESULT_119(RESULT_119),
	.RESULT_120(RESULT_120), .RESULT_121(RESULT_121), .RESULT_122(RESULT_122), .RESULT_123(RESULT_123), .RESULT_124(RESULT_124), .RESULT_125(RESULT_125), .RESULT_126(RESULT_126), .RESULT_127(RESULT_127),
	.RESULT_128(RESULT_128), .RESULT_129(RESULT_129), .RESULT_130(RESULT_130), .RESULT_131(RESULT_131), .RESULT_132(RESULT_132), .RESULT_133(RESULT_133), .RESULT_134(RESULT_134), .RESULT_135(RESULT_135),
	.RESULT_136(RESULT_136), .RESULT_137(RESULT_137), .RESULT_138(RESULT_138), .RESULT_139(RESULT_139), .RESULT_140(RESULT_140), .RESULT_141(RESULT_141), .RESULT_142(RESULT_142), .RESULT_143(RESULT_143),
	.RESULT_144(RESULT_144), .RESULT_145(RESULT_145), .RESULT_146(RESULT_146), .RESULT_147(RESULT_147), .RESULT_148(RESULT_148), .RESULT_149(RESULT_149), .RESULT_150(RESULT_150), .RESULT_151(RESULT_151),
	.RESULT_152(RESULT_152), .RESULT_153(RESULT_153), .RESULT_154(RESULT_154), .RESULT_155(RESULT_155), .RESULT_156(RESULT_156), .RESULT_157(RESULT_157), .RESULT_158(RESULT_158), .RESULT_159(RESULT_159),
	.RESULT_160(RESULT_160), .RESULT_161(RESULT_161), .RESULT_162(RESULT_162), .RESULT_163(RESULT_163), .RESULT_164(RESULT_164), .RESULT_165(RESULT_165), .RESULT_166(RESULT_166), .RESULT_167(RESULT_167),
	.RESULT_168(RESULT_168), .RESULT_169(RESULT_169), .RESULT_170(RESULT_170), .RESULT_171(RESULT_171), .RESULT_172(RESULT_172), .RESULT_173(RESULT_173), .RESULT_174(RESULT_174), .RESULT_175(RESULT_175),
	.RESULT_176(RESULT_176), .RESULT_177(RESULT_177), .RESULT_178(RESULT_178), .RESULT_179(RESULT_179), .RESULT_180(RESULT_180), .RESULT_181(RESULT_181), .RESULT_182(RESULT_182), .RESULT_183(RESULT_183),
	.RESULT_184(RESULT_184), .RESULT_185(RESULT_185), .RESULT_186(RESULT_186), .RESULT_187(RESULT_187), .RESULT_188(RESULT_188), .RESULT_189(RESULT_189), .RESULT_190(RESULT_190), .RESULT_191(RESULT_191),
	.RESULT_192(RESULT_192), .RESULT_193(RESULT_193), .RESULT_194(RESULT_194), .RESULT_195(RESULT_195), .RESULT_196(RESULT_196), .RESULT_197(RESULT_197), .RESULT_198(RESULT_198), .RESULT_199(RESULT_199),
	.RESULT_200(RESULT_200), .RESULT_201(RESULT_201), .RESULT_202(RESULT_202), .RESULT_203(RESULT_203), .RESULT_204(RESULT_204), .RESULT_205(RESULT_205), .RESULT_206(RESULT_206), .RESULT_207(RESULT_207),
	.RESULT_208(RESULT_208), .RESULT_209(RESULT_209), .RESULT_210(RESULT_210), .RESULT_211(RESULT_211), .RESULT_212(RESULT_212), .RESULT_213(RESULT_213), .RESULT_214(RESULT_214), .RESULT_215(RESULT_215),
	.RESULT_216(RESULT_216), .RESULT_217(RESULT_217), .RESULT_218(RESULT_218), .RESULT_219(RESULT_219), .RESULT_220(RESULT_220), .RESULT_221(RESULT_221), .RESULT_222(RESULT_222), .RESULT_223(RESULT_223),
	.RESULT_224(RESULT_224), .RESULT_225(RESULT_225), .RESULT_226(RESULT_226), .RESULT_227(RESULT_227), .RESULT_228(RESULT_228), .RESULT_229(RESULT_229), .RESULT_230(RESULT_230), .RESULT_231(RESULT_231),
	.RESULT_232(RESULT_232), .RESULT_233(RESULT_233), .RESULT_234(RESULT_234), .RESULT_235(RESULT_235), .RESULT_236(RESULT_236), .RESULT_237(RESULT_237), .RESULT_238(RESULT_238), .RESULT_239(RESULT_239),
	.RESULT_240(RESULT_240), .RESULT_241(RESULT_241), .RESULT_242(RESULT_242), .RESULT_243(RESULT_243), .RESULT_244(RESULT_244), .RESULT_245(RESULT_245), .RESULT_246(RESULT_246), .RESULT_247(RESULT_247),
	.RESULT_248(RESULT_248), .RESULT_249(RESULT_249), .RESULT_250(RESULT_250), .RESULT_251(RESULT_251), .RESULT_252(RESULT_252), .RESULT_253(RESULT_253), .RESULT_254(RESULT_254), .RESULT_255(RESULT_255),
	.RESULT_256(RESULT_256), .RESULT_257(RESULT_257), .RESULT_258(RESULT_258), .RESULT_259(RESULT_259), .RESULT_260(RESULT_260), .RESULT_261(RESULT_261), .RESULT_262(RESULT_262), .RESULT_263(RESULT_263),
	.RESULT_264(RESULT_264), .RESULT_265(RESULT_265), .RESULT_266(RESULT_266), .RESULT_267(RESULT_267), .RESULT_268(RESULT_268), .RESULT_269(RESULT_269), .RESULT_270(RESULT_270), .RESULT_271(RESULT_271),
	.RESULT_272(RESULT_272), .RESULT_273(RESULT_273), .RESULT_274(RESULT_274), .RESULT_275(RESULT_275), .RESULT_276(RESULT_276), .RESULT_277(RESULT_277), .RESULT_278(RESULT_278), .RESULT_279(RESULT_279),
	.RESULT_280(RESULT_280), .RESULT_281(RESULT_281), .RESULT_282(RESULT_282), .RESULT_283(RESULT_283), .RESULT_284(RESULT_284), .RESULT_285(RESULT_285), .RESULT_286(RESULT_286), .RESULT_287(RESULT_287),
	.RESULT_288(RESULT_288), .RESULT_289(RESULT_289), .RESULT_290(RESULT_290), .RESULT_291(RESULT_291), .RESULT_292(RESULT_292), .RESULT_293(RESULT_293), .RESULT_294(RESULT_294), .RESULT_295(RESULT_295),
	.RESULT_296(RESULT_296), .RESULT_297(RESULT_297), .RESULT_298(RESULT_298), .RESULT_299(RESULT_299), .RESULT_300(RESULT_300), .RESULT_301(RESULT_301), .RESULT_302(RESULT_302), .RESULT_303(RESULT_303),
	.RESULT_304(RESULT_304), .RESULT_305(RESULT_305), .RESULT_306(RESULT_306), .RESULT_307(RESULT_307), .RESULT_308(RESULT_308), .RESULT_309(RESULT_309), .RESULT_310(RESULT_310), .RESULT_311(RESULT_311),
	.RESULT_312(RESULT_312), .RESULT_313(RESULT_313), .RESULT_314(RESULT_314), .RESULT_315(RESULT_315), .RESULT_316(RESULT_316), .RESULT_317(RESULT_317), .RESULT_318(RESULT_318), .RESULT_319(RESULT_319),
	.RESULT_320(RESULT_320), .RESULT_321(RESULT_321), .RESULT_322(RESULT_322), .RESULT_323(RESULT_323), .RESULT_324(RESULT_324), .RESULT_325(RESULT_325), .RESULT_326(RESULT_326), .RESULT_327(RESULT_327),
	.RESULT_328(RESULT_328), .RESULT_329(RESULT_329), .RESULT_330(RESULT_330), .RESULT_331(RESULT_331), .RESULT_332(RESULT_332), .RESULT_333(RESULT_333), .RESULT_334(RESULT_334), .RESULT_335(RESULT_335),
	.RESULT_336(RESULT_336), .RESULT_337(RESULT_337), .RESULT_338(RESULT_338), .RESULT_339(RESULT_339), .RESULT_340(RESULT_340), .RESULT_341(RESULT_341), .RESULT_342(RESULT_342), .RESULT_343(RESULT_343),
	.RESULT_344(RESULT_344), .RESULT_345(RESULT_345), .RESULT_346(RESULT_346), .RESULT_347(RESULT_347), .RESULT_348(RESULT_348), .RESULT_349(RESULT_349), .RESULT_350(RESULT_350), .RESULT_351(RESULT_351),
	.RESULT_352(RESULT_352), .RESULT_353(RESULT_353), .RESULT_354(RESULT_354), .RESULT_355(RESULT_355), .RESULT_356(RESULT_356), .RESULT_357(RESULT_357), .RESULT_358(RESULT_358), .RESULT_359(RESULT_359),
	.RESULT_360(RESULT_360), .RESULT_361(RESULT_361), .RESULT_362(RESULT_362), .RESULT_363(RESULT_363), .RESULT_364(RESULT_364), .RESULT_365(RESULT_365), .RESULT_366(RESULT_366), .RESULT_367(RESULT_367),
	.RESULT_368(RESULT_368), .RESULT_369(RESULT_369), .RESULT_370(RESULT_370), .RESULT_371(RESULT_371), .RESULT_372(RESULT_372), .RESULT_373(RESULT_373), .RESULT_374(RESULT_374), .RESULT_375(RESULT_375),
	.RESULT_376(RESULT_376), .RESULT_377(RESULT_377), .RESULT_378(RESULT_378), .RESULT_379(RESULT_379), .RESULT_380(RESULT_380), .RESULT_381(RESULT_381), .RESULT_382(RESULT_382), .RESULT_383(RESULT_383),
	.RESULT_384(RESULT_384), .RESULT_385(RESULT_385), .RESULT_386(RESULT_386), .RESULT_387(RESULT_387), .RESULT_388(RESULT_388), .RESULT_389(RESULT_389), .RESULT_390(RESULT_390), .RESULT_391(RESULT_391),
	.RESULT_392(RESULT_392), .RESULT_393(RESULT_393), .RESULT_394(RESULT_394), .RESULT_395(RESULT_395), .RESULT_396(RESULT_396), .RESULT_397(RESULT_397), .RESULT_398(RESULT_398), .RESULT_399(RESULT_399),
	.RESULT_400(RESULT_400), .RESULT_401(RESULT_401), .RESULT_402(RESULT_402), .RESULT_403(RESULT_403), .RESULT_404(RESULT_404), .RESULT_405(RESULT_405), .RESULT_406(RESULT_406), .RESULT_407(RESULT_407),
	.RESULT_408(RESULT_408), .RESULT_409(RESULT_409), .RESULT_410(RESULT_410), .RESULT_411(RESULT_411), .RESULT_412(RESULT_412), .RESULT_413(RESULT_413), .RESULT_414(RESULT_414), .RESULT_415(RESULT_415),
	.RESULT_416(RESULT_416), .RESULT_417(RESULT_417), .RESULT_418(RESULT_418), .RESULT_419(RESULT_419), .RESULT_420(RESULT_420), .RESULT_421(RESULT_421), .RESULT_422(RESULT_422), .RESULT_423(RESULT_423),
	.RESULT_424(RESULT_424), .RESULT_425(RESULT_425), .RESULT_426(RESULT_426), .RESULT_427(RESULT_427), .RESULT_428(RESULT_428), .RESULT_429(RESULT_429), .RESULT_430(RESULT_430), .RESULT_431(RESULT_431),
	.RESULT_432(RESULT_432), .RESULT_433(RESULT_433), .RESULT_434(RESULT_434), .RESULT_435(RESULT_435), .RESULT_436(RESULT_436), .RESULT_437(RESULT_437), .RESULT_438(RESULT_438), .RESULT_439(RESULT_439),
	.RESULT_440(RESULT_440), .RESULT_441(RESULT_441), .RESULT_442(RESULT_442), .RESULT_443(RESULT_443), .RESULT_444(RESULT_444), .RESULT_445(RESULT_445), .RESULT_446(RESULT_446), .RESULT_447(RESULT_447),
	.RESULT_448(RESULT_448), .RESULT_449(RESULT_449), .RESULT_450(RESULT_450), .RESULT_451(RESULT_451), .RESULT_452(RESULT_452), .RESULT_453(RESULT_453), .RESULT_454(RESULT_454), .RESULT_455(RESULT_455),
	.RESULT_456(RESULT_456), .RESULT_457(RESULT_457), .RESULT_458(RESULT_458), .RESULT_459(RESULT_459), .RESULT_460(RESULT_460), .RESULT_461(RESULT_461), .RESULT_462(RESULT_462), .RESULT_463(RESULT_463),
	.RESULT_464(RESULT_464), .RESULT_465(RESULT_465), .RESULT_466(RESULT_466), .RESULT_467(RESULT_467), .RESULT_468(RESULT_468), .RESULT_469(RESULT_469), .RESULT_470(RESULT_470), .RESULT_471(RESULT_471),
	.RESULT_472(RESULT_472), .RESULT_473(RESULT_473), .RESULT_474(RESULT_474), .RESULT_475(RESULT_475), .RESULT_476(RESULT_476), .RESULT_477(RESULT_477), .RESULT_478(RESULT_478), .RESULT_479(RESULT_479),
	.RESULT_480(RESULT_480), .RESULT_481(RESULT_481), .RESULT_482(RESULT_482), .RESULT_483(RESULT_483), .RESULT_484(RESULT_484), .RESULT_485(RESULT_485), .RESULT_486(RESULT_486), .RESULT_487(RESULT_487),
	.RESULT_488(RESULT_488), .RESULT_489(RESULT_489), .RESULT_490(RESULT_490), .RESULT_491(RESULT_491), .RESULT_492(RESULT_492), .RESULT_493(RESULT_493), .RESULT_494(RESULT_494), .RESULT_495(RESULT_495),
	.RESULT_496(RESULT_496), .RESULT_497(RESULT_497), .RESULT_498(RESULT_498), .RESULT_499(RESULT_499), .RESULT_500(RESULT_500), .RESULT_501(RESULT_501), .RESULT_502(RESULT_502), .RESULT_503(RESULT_503),
	.RESULT_504(RESULT_504), .RESULT_505(RESULT_505), .RESULT_506(RESULT_506), .RESULT_507(RESULT_507), .RESULT_508(RESULT_508), .RESULT_509(RESULT_509), .RESULT_510(RESULT_510), .RESULT_511(RESULT_511),
	.RESULT_512(RESULT_512), .RESULT_513(RESULT_513), .RESULT_514(RESULT_514), .RESULT_515(RESULT_515), .RESULT_516(RESULT_516), .RESULT_517(RESULT_517), .RESULT_518(RESULT_518), .RESULT_519(RESULT_519),
	.RESULT_520(RESULT_520), .RESULT_521(RESULT_521), .RESULT_522(RESULT_522), .RESULT_523(RESULT_523), .RESULT_524(RESULT_524), .RESULT_525(RESULT_525), .RESULT_526(RESULT_526), .RESULT_527(RESULT_527),
	.RESULT_528(RESULT_528), .RESULT_529(RESULT_529), .RESULT_530(RESULT_530), .RESULT_531(RESULT_531), .RESULT_532(RESULT_532), .RESULT_533(RESULT_533), .RESULT_534(RESULT_534), .RESULT_535(RESULT_535),
	.RESULT_536(RESULT_536), .RESULT_537(RESULT_537), .RESULT_538(RESULT_538), .RESULT_539(RESULT_539), .RESULT_540(RESULT_540), .RESULT_541(RESULT_541), .RESULT_542(RESULT_542), .RESULT_543(RESULT_543),
	.RESULT_544(RESULT_544), .RESULT_545(RESULT_545), .RESULT_546(RESULT_546), .RESULT_547(RESULT_547), .RESULT_548(RESULT_548), .RESULT_549(RESULT_549), .RESULT_550(RESULT_550), .RESULT_551(RESULT_551),
	.RESULT_552(RESULT_552), .RESULT_553(RESULT_553), .RESULT_554(RESULT_554), .RESULT_555(RESULT_555), .RESULT_556(RESULT_556), .RESULT_557(RESULT_557), .RESULT_558(RESULT_558), .RESULT_559(RESULT_559),
	.RESULT_560(RESULT_560), .RESULT_561(RESULT_561), .RESULT_562(RESULT_562), .RESULT_563(RESULT_563), .RESULT_564(RESULT_564), .RESULT_565(RESULT_565), .RESULT_566(RESULT_566), .RESULT_567(RESULT_567),
	.RESULT_568(RESULT_568), .RESULT_569(RESULT_569), .RESULT_570(RESULT_570), .RESULT_571(RESULT_571), .RESULT_572(RESULT_572), .RESULT_573(RESULT_573), .RESULT_574(RESULT_574), .RESULT_575(RESULT_575),
	.RESULT_576(RESULT_576), .RESULT_577(RESULT_577), .RESULT_578(RESULT_578), .RESULT_579(RESULT_579), .RESULT_580(RESULT_580), .RESULT_581(RESULT_581), .RESULT_582(RESULT_582), .RESULT_583(RESULT_583),
	.RESULT_584(RESULT_584), .RESULT_585(RESULT_585), .RESULT_586(RESULT_586), .RESULT_587(RESULT_587), .RESULT_588(RESULT_588), .RESULT_589(RESULT_589), .RESULT_590(RESULT_590), .RESULT_591(RESULT_591),
	.RESULT_592(RESULT_592), .RESULT_593(RESULT_593), .RESULT_594(RESULT_594), .RESULT_595(RESULT_595), .RESULT_596(RESULT_596), .RESULT_597(RESULT_597), .RESULT_598(RESULT_598), .RESULT_599(RESULT_599),
	.RESULT_600(RESULT_600), .RESULT_601(RESULT_601), .RESULT_602(RESULT_602), .RESULT_603(RESULT_603), .RESULT_604(RESULT_604), .RESULT_605(RESULT_605), .RESULT_606(RESULT_606), .RESULT_607(RESULT_607),
	.RESULT_608(RESULT_608), .RESULT_609(RESULT_609), .RESULT_610(RESULT_610), .RESULT_611(RESULT_611), .RESULT_612(RESULT_612), .RESULT_613(RESULT_613), .RESULT_614(RESULT_614), .RESULT_615(RESULT_615),
	.RESULT_616(RESULT_616), .RESULT_617(RESULT_617), .RESULT_618(RESULT_618), .RESULT_619(RESULT_619), .RESULT_620(RESULT_620), .RESULT_621(RESULT_621), .RESULT_622(RESULT_622), .RESULT_623(RESULT_623),
	.RESULT_624(RESULT_624), .RESULT_625(RESULT_625), .RESULT_626(RESULT_626), .RESULT_627(RESULT_627), .RESULT_628(RESULT_628), .RESULT_629(RESULT_629), .RESULT_630(RESULT_630), .RESULT_631(RESULT_631),
	.RESULT_632(RESULT_632), .RESULT_633(RESULT_633), .RESULT_634(RESULT_634), .RESULT_635(RESULT_635), .RESULT_636(RESULT_636), .RESULT_637(RESULT_637), .RESULT_638(RESULT_638), .RESULT_639(RESULT_639),
	.RESULT_640(RESULT_640), .RESULT_641(RESULT_641), .RESULT_642(RESULT_642), .RESULT_643(RESULT_643), .RESULT_644(RESULT_644), .RESULT_645(RESULT_645), .RESULT_646(RESULT_646), .RESULT_647(RESULT_647),
	.RESULT_648(RESULT_648), .RESULT_649(RESULT_649), .RESULT_650(RESULT_650), .RESULT_651(RESULT_651), .RESULT_652(RESULT_652), .RESULT_653(RESULT_653), .RESULT_654(RESULT_654), .RESULT_655(RESULT_655),
	.RESULT_656(RESULT_656), .RESULT_657(RESULT_657), .RESULT_658(RESULT_658), .RESULT_659(RESULT_659), .RESULT_660(RESULT_660), .RESULT_661(RESULT_661), .RESULT_662(RESULT_662), .RESULT_663(RESULT_663),
	.RESULT_664(RESULT_664), .RESULT_665(RESULT_665), .RESULT_666(RESULT_666), .RESULT_667(RESULT_667), .RESULT_668(RESULT_668), .RESULT_669(RESULT_669), .RESULT_670(RESULT_670), .RESULT_671(RESULT_671),
	.RESULT_672(RESULT_672), .RESULT_673(RESULT_673), .RESULT_674(RESULT_674), .RESULT_675(RESULT_675), .RESULT_676(RESULT_676), .RESULT_677(RESULT_677), .RESULT_678(RESULT_678), .RESULT_679(RESULT_679),
	.RESULT_680(RESULT_680), .RESULT_681(RESULT_681), .RESULT_682(RESULT_682), .RESULT_683(RESULT_683),
	.RESULT_684(RESULT_684), .RESULT_685(RESULT_685), .RESULT_686(RESULT_686), .RESULT_687(RESULT_687),
	.RESULT_688(RESULT_688), .RESULT_689(RESULT_689), .RESULT_690(RESULT_690), .RESULT_691(RESULT_691),
	.RESULT_692(RESULT_692), .RESULT_693(RESULT_693), .RESULT_694(RESULT_694), .RESULT_695(RESULT_695),
	.RESULT_696(RESULT_696), .RESULT_697(RESULT_697), .RESULT_698(RESULT_698), .RESULT_699(RESULT_699),
	.RESULT_700(RESULT_700), .RESULT_701(RESULT_701), .RESULT_702(RESULT_702), .RESULT_703(RESULT_703),
	.RESULT_704(RESULT_704), .RESULT_705(RESULT_705), .RESULT_706(RESULT_706), .RESULT_707(RESULT_707),
	.RESULT_708(RESULT_708), .RESULT_709(RESULT_709), .RESULT_710(RESULT_710), .RESULT_711(RESULT_711),
	.RESULT_712(RESULT_712), .RESULT_713(RESULT_713), .RESULT_714(RESULT_714), .RESULT_715(RESULT_715),
	.RESULT_716(RESULT_716), .RESULT_717(RESULT_717), .RESULT_718(RESULT_718), .RESULT_719(RESULT_719),
	.RESULT_720(RESULT_720), .RESULT_721(RESULT_721), .RESULT_722(RESULT_722), .RESULT_723(RESULT_723),
	.RESULT_724(RESULT_724), .RESULT_725(RESULT_725), .RESULT_726(RESULT_726), .RESULT_727(RESULT_727),
	.RESULT_728(RESULT_728), .RESULT_729(RESULT_729), .RESULT_730(RESULT_730), .RESULT_731(RESULT_731),
	.RESULT_732(RESULT_732), .RESULT_733(RESULT_733), .RESULT_734(RESULT_734), .RESULT_735(RESULT_735),
	.RESULT_736(RESULT_736), .RESULT_737(RESULT_737), .RESULT_738(RESULT_738), .RESULT_739(RESULT_739),
	.RESULT_740(RESULT_740), .RESULT_741(RESULT_741), .RESULT_742(RESULT_742), .RESULT_743(RESULT_743),
	.RESULT_744(RESULT_744), .RESULT_745(RESULT_745), .RESULT_746(RESULT_746), .RESULT_747(RESULT_747),
	.RESULT_748(RESULT_748), .RESULT_749(RESULT_749), .RESULT_750(RESULT_750), .RESULT_751(RESULT_751),
	.RESULT_752(RESULT_752), .RESULT_753(RESULT_753), .RESULT_754(RESULT_754), .RESULT_755(RESULT_755),
	.RESULT_756(RESULT_756), .RESULT_757(RESULT_757), .RESULT_758(RESULT_758), .RESULT_759(RESULT_759),
	.RESULT_760(RESULT_760), .RESULT_761(RESULT_761), .RESULT_762(RESULT_762), .RESULT_763(RESULT_763),
	.RESULT_764(RESULT_764), .RESULT_765(RESULT_765), .RESULT_766(RESULT_766), .RESULT_767(RESULT_767),
	.RESULT_768(RESULT_768), .RESULT_769(RESULT_769), .RESULT_770(RESULT_770), .RESULT_771(RESULT_771),
	.RESULT_772(RESULT_772), .RESULT_773(RESULT_773), .RESULT_774(RESULT_774), .RESULT_775(RESULT_775),
	.RESULT_776(RESULT_776), .RESULT_777(RESULT_777), .RESULT_778(RESULT_778), .RESULT_779(RESULT_779),
	.RESULT_780(RESULT_780), .RESULT_781(RESULT_781), .RESULT_782(RESULT_782), .RESULT_783(RESULT_783),
	.RESULT_784(RESULT_784), .RESULT_785(RESULT_785), .RESULT_786(RESULT_786), .RESULT_787(RESULT_787),
	.RESULT_788(RESULT_788), .RESULT_789(RESULT_789), .RESULT_790(RESULT_790), .RESULT_791(RESULT_791),
	.RESULT_792(RESULT_792), .RESULT_793(RESULT_793), .RESULT_794(RESULT_794), .RESULT_795(RESULT_795),
	.RESULT_796(RESULT_796), .RESULT_797(RESULT_797), .RESULT_798(RESULT_798), .RESULT_799(RESULT_799),
	.RESULT_800(RESULT_800), .RESULT_801(RESULT_801), .RESULT_802(RESULT_802), .RESULT_803(RESULT_803),
	.RESULT_804(RESULT_804), .RESULT_805(RESULT_805), .RESULT_806(RESULT_806), .RESULT_807(RESULT_807),
	.RESULT_808(RESULT_808), .RESULT_809(RESULT_809), .RESULT_810(RESULT_810), .RESULT_811(RESULT_811),
	.RESULT_812(RESULT_812), .RESULT_813(RESULT_813), .RESULT_814(RESULT_814), .RESULT_815(RESULT_815),
	.RESULT_816(RESULT_816), .RESULT_817(RESULT_817), .RESULT_818(RESULT_818), .RESULT_819(RESULT_819),
	.RESULT_820(RESULT_820), .RESULT_821(RESULT_821), .RESULT_822(RESULT_822), .RESULT_823(RESULT_823),
	.RESULT_824(RESULT_824), .RESULT_825(RESULT_825), .RESULT_826(RESULT_826), .RESULT_827(RESULT_827),
	.RESULT_828(RESULT_828), .RESULT_829(RESULT_829), .RESULT_830(RESULT_830), .RESULT_831(RESULT_831),
	.RESULT_832(RESULT_832), .RESULT_833(RESULT_833), .RESULT_834(RESULT_834), .RESULT_835(RESULT_835),
	.RESULT_836(RESULT_836), .RESULT_837(RESULT_837), .RESULT_838(RESULT_838), .RESULT_839(RESULT_839),
	.RESULT_840(RESULT_840), .RESULT_841(RESULT_841), .RESULT_842(RESULT_842), .RESULT_843(RESULT_843),
	.RESULT_844(RESULT_844), .RESULT_845(RESULT_845), .RESULT_846(RESULT_846), .RESULT_847(RESULT_847),
	.RESULT_848(RESULT_848), .RESULT_849(RESULT_849), .RESULT_850(RESULT_850), .RESULT_851(RESULT_851),
	.RESULT_852(RESULT_852), .RESULT_853(RESULT_853), .RESULT_854(RESULT_854), .RESULT_855(RESULT_855),
	.RESULT_856(RESULT_856), .RESULT_857(RESULT_857), .RESULT_858(RESULT_858), .RESULT_859(RESULT_859),
	.RESULT_860(RESULT_860), .RESULT_861(RESULT_861), .RESULT_862(RESULT_862), .RESULT_863(RESULT_863),
	.RESULT_864(RESULT_864), .RESULT_865(RESULT_865), .RESULT_866(RESULT_866), .RESULT_867(RESULT_867),
	.RESULT_868(RESULT_868), .RESULT_869(RESULT_869), .RESULT_870(RESULT_870), .RESULT_871(RESULT_871),
	.RESULT_872(RESULT_872), .RESULT_873(RESULT_873), .RESULT_874(RESULT_874), .RESULT_875(RESULT_875),
	.RESULT_876(RESULT_876), .RESULT_877(RESULT_877), .RESULT_878(RESULT_878), .RESULT_879(RESULT_879),
	.RESULT_880(RESULT_880), .RESULT_881(RESULT_881), .RESULT_882(RESULT_882), .RESULT_883(RESULT_883),
	.RESULT_884(RESULT_884), .RESULT_885(RESULT_885), .RESULT_886(RESULT_886), .RESULT_887(RESULT_887),
	.RESULT_888(RESULT_888), .RESULT_889(RESULT_889), .RESULT_890(RESULT_890), .RESULT_891(RESULT_891),
	.RESULT_892(RESULT_892), .RESULT_893(RESULT_893), .RESULT_894(RESULT_894), .RESULT_895(RESULT_895)
);
endmodule
