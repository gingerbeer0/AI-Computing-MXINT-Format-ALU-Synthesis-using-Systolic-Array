module output_buffer(
   input CLK,
   input RSTN,
   input result_enable,
   input signed [15:0] RESULT_P18, // Output array
   input signed [15:0] RESULT_P17, // Output array
   input signed [15:0] RESULT_P16, // Output array
   input signed [15:0] RESULT_P15, // Output array
   input signed [15:0] RESULT_P14, // Output array
   input signed [15:0] RESULT_P13, // Output array
   input signed [15:0] RESULT_P12, // Output array
   input signed [15:0] RESULT_P28, // Output array
   input signed [15:0] RESULT_P27, // Output array
   input signed [15:0] RESULT_P26, // Output array
   input signed [15:0] RESULT_P25, // Output array
   input signed [15:0] RESULT_P24, // Output array
   input signed [15:0] RESULT_P23, // Output array
   input signed [15:0] RESULT_P38, // Output array
   input signed [15:0] RESULT_P37, // Output array
   input signed [15:0] RESULT_P36, // Output array
   input signed [15:0] RESULT_P35, // Output array
   input signed [15:0] RESULT_P34, // Output array
   input signed [15:0] RESULT_P48, // Output array
   input signed [15:0] RESULT_P47, // Output array
   input signed [15:0] RESULT_P46, // Output array
   input signed [15:0] RESULT_P45, // Output array
   input signed [15:0] RESULT_P58, // Output array
   input signed [15:0] RESULT_P57, // Output array
   input signed [15:0] RESULT_P56, // Output array
   input signed [15:0] RESULT_P68, // Output array
   input signed [15:0] RESULT_P67, // Output array
   input signed [15:0] RESULT_P78, // Output array

   output reg signed [15:0] RESULT_0,
output reg signed [15:0] RESULT_1,
output reg signed [15:0] RESULT_2,
output reg signed [15:0] RESULT_3,
output reg signed [15:0] RESULT_4,
output reg signed [15:0] RESULT_5,
output reg signed [15:0] RESULT_6,
output reg signed [15:0] RESULT_7,
output reg signed [15:0] RESULT_8,
output reg signed [15:0] RESULT_9,
output reg signed [15:0] RESULT_10,
output reg signed [15:0] RESULT_11,
output reg signed [15:0] RESULT_12,
output reg signed [15:0] RESULT_13,
output reg signed [15:0] RESULT_14,
output reg signed [15:0] RESULT_15,
output reg signed [15:0] RESULT_16,
output reg signed [15:0] RESULT_17,
output reg signed [15:0] RESULT_18,
output reg signed [15:0] RESULT_19,
output reg signed [15:0] RESULT_20,
output reg signed [15:0] RESULT_21,
output reg signed [15:0] RESULT_22,
output reg signed [15:0] RESULT_23,
output reg signed [15:0] RESULT_24,
output reg signed [15:0] RESULT_25,
output reg signed [15:0] RESULT_26,
output reg signed [15:0] RESULT_27,
output reg signed [15:0] RESULT_28,
output reg signed [15:0] RESULT_29,
output reg signed [15:0] RESULT_30,
output reg signed [15:0] RESULT_31,
output reg signed [15:0] RESULT_32,
output reg signed [15:0] RESULT_33,
output reg signed [15:0] RESULT_34,
output reg signed [15:0] RESULT_35,
output reg signed [15:0] RESULT_36,
output reg signed [15:0] RESULT_37,
output reg signed [15:0] RESULT_38,
output reg signed [15:0] RESULT_39,
output reg signed [15:0] RESULT_40,
output reg signed [15:0] RESULT_41,
output reg signed [15:0] RESULT_42,
output reg signed [15:0] RESULT_43,
output reg signed [15:0] RESULT_44,
output reg signed [15:0] RESULT_45,
output reg signed [15:0] RESULT_46,
output reg signed [15:0] RESULT_47,
output reg signed [15:0] RESULT_48,
output reg signed [15:0] RESULT_49,
output reg signed [15:0] RESULT_50,
output reg signed [15:0] RESULT_51,
output reg signed [15:0] RESULT_52,
output reg signed [15:0] RESULT_53,
output reg signed [15:0] RESULT_54,
output reg signed [15:0] RESULT_55,
output reg signed [15:0] RESULT_56,
output reg signed [15:0] RESULT_57,
output reg signed [15:0] RESULT_58,
output reg signed [15:0] RESULT_59,
output reg signed [15:0] RESULT_60,
output reg signed [15:0] RESULT_61,
output reg signed [15:0] RESULT_62,
output reg signed [15:0] RESULT_63,
output reg signed [15:0] RESULT_64,
output reg signed [15:0] RESULT_65,
output reg signed [15:0] RESULT_66,
output reg signed [15:0] RESULT_67,
output reg signed [15:0] RESULT_68,
output reg signed [15:0] RESULT_69,
output reg signed [15:0] RESULT_70,
output reg signed [15:0] RESULT_71,
output reg signed [15:0] RESULT_72,
output reg signed [15:0] RESULT_73,
output reg signed [15:0] RESULT_74,
output reg signed [15:0] RESULT_75,
output reg signed [15:0] RESULT_76,
output reg signed [15:0] RESULT_77,
output reg signed [15:0] RESULT_78,
output reg signed [15:0] RESULT_79,
output reg signed [15:0] RESULT_80,
output reg signed [15:0] RESULT_81,
output reg signed [15:0] RESULT_82,
output reg signed [15:0] RESULT_83,
output reg signed [15:0] RESULT_84,
output reg signed [15:0] RESULT_85,
output reg signed [15:0] RESULT_86,
output reg signed [15:0] RESULT_87,
output reg signed [15:0] RESULT_88,
output reg signed [15:0] RESULT_89,
output reg signed [15:0] RESULT_90,
output reg signed [15:0] RESULT_91,
output reg signed [15:0] RESULT_92,
output reg signed [15:0] RESULT_93,
output reg signed [15:0] RESULT_94,
output reg signed [15:0] RESULT_95,
output reg signed [15:0] RESULT_96,
output reg signed [15:0] RESULT_97,
output reg signed [15:0] RESULT_98,
output reg signed [15:0] RESULT_99,
output reg signed [15:0] RESULT_100,
output reg signed [15:0] RESULT_101,
output reg signed [15:0] RESULT_102,
output reg signed [15:0] RESULT_103,
output reg signed [15:0] RESULT_104,
output reg signed [15:0] RESULT_105,
output reg signed [15:0] RESULT_106,
output reg signed [15:0] RESULT_107,
output reg signed [15:0] RESULT_108,
output reg signed [15:0] RESULT_109,
output reg signed [15:0] RESULT_110,
output reg signed [15:0] RESULT_111,
output reg signed [15:0] RESULT_112,
output reg signed [15:0] RESULT_113,
output reg signed [15:0] RESULT_114,
output reg signed [15:0] RESULT_115,
output reg signed [15:0] RESULT_116,
output reg signed [15:0] RESULT_117,
output reg signed [15:0] RESULT_118,
output reg signed [15:0] RESULT_119,
output reg signed [15:0] RESULT_120,
output reg signed [15:0] RESULT_121,
output reg signed [15:0] RESULT_122,
output reg signed [15:0] RESULT_123,
output reg signed [15:0] RESULT_124,
output reg signed [15:0] RESULT_125,
output reg signed [15:0] RESULT_126,
output reg signed [15:0] RESULT_127,
output reg signed [15:0] RESULT_128,
output reg signed [15:0] RESULT_129,
output reg signed [15:0] RESULT_130,
output reg signed [15:0] RESULT_131,
output reg signed [15:0] RESULT_132,
output reg signed [15:0] RESULT_133,
output reg signed [15:0] RESULT_134,
output reg signed [15:0] RESULT_135,
output reg signed [15:0] RESULT_136,
output reg signed [15:0] RESULT_137,
output reg signed [15:0] RESULT_138,
output reg signed [15:0] RESULT_139,
output reg signed [15:0] RESULT_140,
output reg signed [15:0] RESULT_141,
output reg signed [15:0] RESULT_142,
output reg signed [15:0] RESULT_143,
output reg signed [15:0] RESULT_144,
output reg signed [15:0] RESULT_145,
output reg signed [15:0] RESULT_146,
output reg signed [15:0] RESULT_147,
output reg signed [15:0] RESULT_148,
output reg signed [15:0] RESULT_149,
output reg signed [15:0] RESULT_150,
output reg signed [15:0] RESULT_151,
output reg signed [15:0] RESULT_152,
output reg signed [15:0] RESULT_153,
output reg signed [15:0] RESULT_154,
output reg signed [15:0] RESULT_155,
output reg signed [15:0] RESULT_156,
output reg signed [15:0] RESULT_157,
output reg signed [15:0] RESULT_158,
output reg signed [15:0] RESULT_159,
output reg signed [15:0] RESULT_160,
output reg signed [15:0] RESULT_161,
output reg signed [15:0] RESULT_162,
output reg signed [15:0] RESULT_163,
output reg signed [15:0] RESULT_164,
output reg signed [15:0] RESULT_165,
output reg signed [15:0] RESULT_166,
output reg signed [15:0] RESULT_167,
output reg signed [15:0] RESULT_168,
output reg signed [15:0] RESULT_169,
output reg signed [15:0] RESULT_170,
output reg signed [15:0] RESULT_171,
output reg signed [15:0] RESULT_172,
output reg signed [15:0] RESULT_173,
output reg signed [15:0] RESULT_174,
output reg signed [15:0] RESULT_175,
output reg signed [15:0] RESULT_176,
output reg signed [15:0] RESULT_177,
output reg signed [15:0] RESULT_178,
output reg signed [15:0] RESULT_179,
output reg signed [15:0] RESULT_180,
output reg signed [15:0] RESULT_181,
output reg signed [15:0] RESULT_182,
output reg signed [15:0] RESULT_183,
output reg signed [15:0] RESULT_184,
output reg signed [15:0] RESULT_185,
output reg signed [15:0] RESULT_186,
output reg signed [15:0] RESULT_187,
output reg signed [15:0] RESULT_188,
output reg signed [15:0] RESULT_189,
output reg signed [15:0] RESULT_190,
output reg signed [15:0] RESULT_191,
output reg signed [15:0] RESULT_192,
output reg signed [15:0] RESULT_193,
output reg signed [15:0] RESULT_194,
output reg signed [15:0] RESULT_195,
output reg signed [15:0] RESULT_196,
output reg signed [15:0] RESULT_197,
output reg signed [15:0] RESULT_198,
output reg signed [15:0] RESULT_199,
output reg signed [15:0] RESULT_200,
output reg signed [15:0] RESULT_201,
output reg signed [15:0] RESULT_202,
output reg signed [15:0] RESULT_203,
output reg signed [15:0] RESULT_204,
output reg signed [15:0] RESULT_205,
output reg signed [15:0] RESULT_206,
output reg signed [15:0] RESULT_207,
output reg signed [15:0] RESULT_208,
output reg signed [15:0] RESULT_209,
output reg signed [15:0] RESULT_210,
output reg signed [15:0] RESULT_211,
output reg signed [15:0] RESULT_212,
output reg signed [15:0] RESULT_213,
output reg signed [15:0] RESULT_214,
output reg signed [15:0] RESULT_215,
output reg signed [15:0] RESULT_216,
output reg signed [15:0] RESULT_217,
output reg signed [15:0] RESULT_218,
output reg signed [15:0] RESULT_219,
output reg signed [15:0] RESULT_220,
output reg signed [15:0] RESULT_221,
output reg signed [15:0] RESULT_222,
output reg signed [15:0] RESULT_223,
output reg signed [15:0] RESULT_224,
output reg signed [15:0] RESULT_225,
output reg signed [15:0] RESULT_226,
output reg signed [15:0] RESULT_227,
output reg signed [15:0] RESULT_228,
output reg signed [15:0] RESULT_229,
output reg signed [15:0] RESULT_230,
output reg signed [15:0] RESULT_231,
output reg signed [15:0] RESULT_232,
output reg signed [15:0] RESULT_233,
output reg signed [15:0] RESULT_234,
output reg signed [15:0] RESULT_235,
output reg signed [15:0] RESULT_236,
output reg signed [15:0] RESULT_237,
output reg signed [15:0] RESULT_238,
output reg signed [15:0] RESULT_239,
output reg signed [15:0] RESULT_240,
output reg signed [15:0] RESULT_241,
output reg signed [15:0] RESULT_242,
output reg signed [15:0] RESULT_243,
output reg signed [15:0] RESULT_244,
output reg signed [15:0] RESULT_245,
output reg signed [15:0] RESULT_246,
output reg signed [15:0] RESULT_247,
output reg signed [15:0] RESULT_248,
output reg signed [15:0] RESULT_249,
output reg signed [15:0] RESULT_250,
output reg signed [15:0] RESULT_251,
output reg signed [15:0] RESULT_252,
output reg signed [15:0] RESULT_253,
output reg signed [15:0] RESULT_254,
output reg signed [15:0] RESULT_255,
output reg signed [15:0] RESULT_256,
output reg signed [15:0] RESULT_257,
output reg signed [15:0] RESULT_258,
output reg signed [15:0] RESULT_259,
output reg signed [15:0] RESULT_260,
output reg signed [15:0] RESULT_261,
output reg signed [15:0] RESULT_262,
output reg signed [15:0] RESULT_263,
output reg signed [15:0] RESULT_264,
output reg signed [15:0] RESULT_265,
output reg signed [15:0] RESULT_266,
output reg signed [15:0] RESULT_267,
output reg signed [15:0] RESULT_268,
output reg signed [15:0] RESULT_269,
output reg signed [15:0] RESULT_270,
output reg signed [15:0] RESULT_271,
output reg signed [15:0] RESULT_272,
output reg signed [15:0] RESULT_273,
output reg signed [15:0] RESULT_274,
output reg signed [15:0] RESULT_275,
output reg signed [15:0] RESULT_276,
output reg signed [15:0] RESULT_277,
output reg signed [15:0] RESULT_278,
output reg signed [15:0] RESULT_279,
output reg signed [15:0] RESULT_280,
output reg signed [15:0] RESULT_281,
output reg signed [15:0] RESULT_282,
output reg signed [15:0] RESULT_283,
output reg signed [15:0] RESULT_284,
output reg signed [15:0] RESULT_285,
output reg signed [15:0] RESULT_286,
output reg signed [15:0] RESULT_287,
output reg signed [15:0] RESULT_288,
output reg signed [15:0] RESULT_289,
output reg signed [15:0] RESULT_290,
output reg signed [15:0] RESULT_291,
output reg signed [15:0] RESULT_292,
output reg signed [15:0] RESULT_293,
output reg signed [15:0] RESULT_294,
output reg signed [15:0] RESULT_295,
output reg signed [15:0] RESULT_296,
output reg signed [15:0] RESULT_297,
output reg signed [15:0] RESULT_298,
output reg signed [15:0] RESULT_299,
output reg signed [15:0] RESULT_300,
output reg signed [15:0] RESULT_301,
output reg signed [15:0] RESULT_302,
output reg signed [15:0] RESULT_303,
output reg signed [15:0] RESULT_304,
output reg signed [15:0] RESULT_305,
output reg signed [15:0] RESULT_306,
output reg signed [15:0] RESULT_307,
output reg signed [15:0] RESULT_308,
output reg signed [15:0] RESULT_309,
output reg signed [15:0] RESULT_310,
output reg signed [15:0] RESULT_311,
output reg signed [15:0] RESULT_312,
output reg signed [15:0] RESULT_313,
output reg signed [15:0] RESULT_314,
output reg signed [15:0] RESULT_315,
output reg signed [15:0] RESULT_316,
output reg signed [15:0] RESULT_317,
output reg signed [15:0] RESULT_318,
output reg signed [15:0] RESULT_319,
output reg signed [15:0] RESULT_320,
output reg signed [15:0] RESULT_321,
output reg signed [15:0] RESULT_322,
output reg signed [15:0] RESULT_323,
output reg signed [15:0] RESULT_324,
output reg signed [15:0] RESULT_325,
output reg signed [15:0] RESULT_326,
output reg signed [15:0] RESULT_327,
output reg signed [15:0] RESULT_328,
output reg signed [15:0] RESULT_329,
output reg signed [15:0] RESULT_330,
output reg signed [15:0] RESULT_331,
output reg signed [15:0] RESULT_332,
output reg signed [15:0] RESULT_333,
output reg signed [15:0] RESULT_334,
output reg signed [15:0] RESULT_335,
output reg signed [15:0] RESULT_336,
output reg signed [15:0] RESULT_337,
output reg signed [15:0] RESULT_338,
output reg signed [15:0] RESULT_339,
output reg signed [15:0] RESULT_340,
output reg signed [15:0] RESULT_341,
output reg signed [15:0] RESULT_342,
output reg signed [15:0] RESULT_343,
output reg signed [15:0] RESULT_344,
output reg signed [15:0] RESULT_345,
output reg signed [15:0] RESULT_346,
output reg signed [15:0] RESULT_347,
output reg signed [15:0] RESULT_348,
output reg signed [15:0] RESULT_349,
output reg signed [15:0] RESULT_350,
output reg signed [15:0] RESULT_351,
output reg signed [15:0] RESULT_352,
output reg signed [15:0] RESULT_353,
output reg signed [15:0] RESULT_354,
output reg signed [15:0] RESULT_355,
output reg signed [15:0] RESULT_356,
output reg signed [15:0] RESULT_357,
output reg signed [15:0] RESULT_358,
output reg signed [15:0] RESULT_359,
output reg signed [15:0] RESULT_360,
output reg signed [15:0] RESULT_361,
output reg signed [15:0] RESULT_362,
output reg signed [15:0] RESULT_363,
output reg signed [15:0] RESULT_364,
output reg signed [15:0] RESULT_365,
output reg signed [15:0] RESULT_366,
output reg signed [15:0] RESULT_367,
output reg signed [15:0] RESULT_368,
output reg signed [15:0] RESULT_369,
output reg signed [15:0] RESULT_370,
output reg signed [15:0] RESULT_371,
output reg signed [15:0] RESULT_372,
output reg signed [15:0] RESULT_373,
output reg signed [15:0] RESULT_374,
output reg signed [15:0] RESULT_375,
output reg signed [15:0] RESULT_376,
output reg signed [15:0] RESULT_377,
output reg signed [15:0] RESULT_378,
output reg signed [15:0] RESULT_379,
output reg signed [15:0] RESULT_380,
output reg signed [15:0] RESULT_381,
output reg signed [15:0] RESULT_382,
output reg signed [15:0] RESULT_383,
output reg signed [15:0] RESULT_384,
output reg signed [15:0] RESULT_385,
output reg signed [15:0] RESULT_386,
output reg signed [15:0] RESULT_387,
output reg signed [15:0] RESULT_388,
output reg signed [15:0] RESULT_389,
output reg signed [15:0] RESULT_390,
output reg signed [15:0] RESULT_391,
output reg signed [15:0] RESULT_392,
output reg signed [15:0] RESULT_393,
output reg signed [15:0] RESULT_394,
output reg signed [15:0] RESULT_395,
output reg signed [15:0] RESULT_396,
output reg signed [15:0] RESULT_397,
output reg signed [15:0] RESULT_398,
output reg signed [15:0] RESULT_399,
output reg signed [15:0] RESULT_400,
output reg signed [15:0] RESULT_401,
output reg signed [15:0] RESULT_402,
output reg signed [15:0] RESULT_403,
output reg signed [15:0] RESULT_404,
output reg signed [15:0] RESULT_405,
output reg signed [15:0] RESULT_406,
output reg signed [15:0] RESULT_407,
output reg signed [15:0] RESULT_408,
output reg signed [15:0] RESULT_409,
output reg signed [15:0] RESULT_410,
output reg signed [15:0] RESULT_411,
output reg signed [15:0] RESULT_412,
output reg signed [15:0] RESULT_413,
output reg signed [15:0] RESULT_414,
output reg signed [15:0] RESULT_415,
output reg signed [15:0] RESULT_416,
output reg signed [15:0] RESULT_417,
output reg signed [15:0] RESULT_418,
output reg signed [15:0] RESULT_419,
output reg signed [15:0] RESULT_420,
output reg signed [15:0] RESULT_421,
output reg signed [15:0] RESULT_422,
output reg signed [15:0] RESULT_423,
output reg signed [15:0] RESULT_424,
output reg signed [15:0] RESULT_425,
output reg signed [15:0] RESULT_426,
output reg signed [15:0] RESULT_427,
output reg signed [15:0] RESULT_428,
output reg signed [15:0] RESULT_429,
output reg signed [15:0] RESULT_430,
output reg signed [15:0] RESULT_431,
output reg signed [15:0] RESULT_432,
output reg signed [15:0] RESULT_433,
output reg signed [15:0] RESULT_434,
output reg signed [15:0] RESULT_435,
output reg signed [15:0] RESULT_436,
output reg signed [15:0] RESULT_437,
output reg signed [15:0] RESULT_438,
output reg signed [15:0] RESULT_439,
output reg signed [15:0] RESULT_440,
output reg signed [15:0] RESULT_441,
output reg signed [15:0] RESULT_442,
output reg signed [15:0] RESULT_443,
output reg signed [15:0] RESULT_444,
output reg signed [15:0] RESULT_445,
output reg signed [15:0] RESULT_446,
output reg signed [15:0] RESULT_447,
output reg signed [15:0] RESULT_448,
output reg signed [15:0] RESULT_449,
output reg signed [15:0] RESULT_450,
output reg signed [15:0] RESULT_451,
output reg signed [15:0] RESULT_452,
output reg signed [15:0] RESULT_453,
output reg signed [15:0] RESULT_454,
output reg signed [15:0] RESULT_455,
output reg signed [15:0] RESULT_456,
output reg signed [15:0] RESULT_457,
output reg signed [15:0] RESULT_458,
output reg signed [15:0] RESULT_459,
output reg signed [15:0] RESULT_460,
output reg signed [15:0] RESULT_461,
output reg signed [15:0] RESULT_462,
output reg signed [15:0] RESULT_463,
output reg signed [15:0] RESULT_464,
output reg signed [15:0] RESULT_465,
output reg signed [15:0] RESULT_466,
output reg signed [15:0] RESULT_467,
output reg signed [15:0] RESULT_468,
output reg signed [15:0] RESULT_469,
output reg signed [15:0] RESULT_470,
output reg signed [15:0] RESULT_471,
output reg signed [15:0] RESULT_472,
output reg signed [15:0] RESULT_473,
output reg signed [15:0] RESULT_474,
output reg signed [15:0] RESULT_475,
output reg signed [15:0] RESULT_476,
output reg signed [15:0] RESULT_477,
output reg signed [15:0] RESULT_478,
output reg signed [15:0] RESULT_479,
output reg signed [15:0] RESULT_480,
output reg signed [15:0] RESULT_481,
output reg signed [15:0] RESULT_482,
output reg signed [15:0] RESULT_483,
output reg signed [15:0] RESULT_484,
output reg signed [15:0] RESULT_485,
output reg signed [15:0] RESULT_486,
output reg signed [15:0] RESULT_487,
output reg signed [15:0] RESULT_488,
output reg signed [15:0] RESULT_489,
output reg signed [15:0] RESULT_490,
output reg signed [15:0] RESULT_491,
output reg signed [15:0] RESULT_492,
output reg signed [15:0] RESULT_493,
output reg signed [15:0] RESULT_494,
output reg signed [15:0] RESULT_495,
output reg signed [15:0] RESULT_496,
output reg signed [15:0] RESULT_497,
output reg signed [15:0] RESULT_498,
output reg signed [15:0] RESULT_499,
output reg signed [15:0] RESULT_500,
output reg signed [15:0] RESULT_501,
output reg signed [15:0] RESULT_502,
output reg signed [15:0] RESULT_503,
output reg signed [15:0] RESULT_504,
output reg signed [15:0] RESULT_505,
output reg signed [15:0] RESULT_506,
output reg signed [15:0] RESULT_507,
output reg signed [15:0] RESULT_508,
output reg signed [15:0] RESULT_509,
output reg signed [15:0] RESULT_510,
output reg signed [15:0] RESULT_511,
output reg signed [15:0] RESULT_512,
output reg signed [15:0] RESULT_513,
output reg signed [15:0] RESULT_514,
output reg signed [15:0] RESULT_515,
output reg signed [15:0] RESULT_516,
output reg signed [15:0] RESULT_517,
output reg signed [15:0] RESULT_518,
output reg signed [15:0] RESULT_519,
output reg signed [15:0] RESULT_520,
output reg signed [15:0] RESULT_521,
output reg signed [15:0] RESULT_522,
output reg signed [15:0] RESULT_523,
output reg signed [15:0] RESULT_524,
output reg signed [15:0] RESULT_525,
output reg signed [15:0] RESULT_526,
output reg signed [15:0] RESULT_527,
output reg signed [15:0] RESULT_528,
output reg signed [15:0] RESULT_529,
output reg signed [15:0] RESULT_530,
output reg signed [15:0] RESULT_531,
output reg signed [15:0] RESULT_532,
output reg signed [15:0] RESULT_533,
output reg signed [15:0] RESULT_534,
output reg signed [15:0] RESULT_535,
output reg signed [15:0] RESULT_536,
output reg signed [15:0] RESULT_537,
output reg signed [15:0] RESULT_538,
output reg signed [15:0] RESULT_539,
output reg signed [15:0] RESULT_540,
output reg signed [15:0] RESULT_541,
output reg signed [15:0] RESULT_542,
output reg signed [15:0] RESULT_543,
output reg signed [15:0] RESULT_544,
output reg signed [15:0] RESULT_545,
output reg signed [15:0] RESULT_546,
output reg signed [15:0] RESULT_547,
output reg signed [15:0] RESULT_548,
output reg signed [15:0] RESULT_549,
output reg signed [15:0] RESULT_550,
output reg signed [15:0] RESULT_551,
output reg signed [15:0] RESULT_552,
output reg signed [15:0] RESULT_553,
output reg signed [15:0] RESULT_554,
output reg signed [15:0] RESULT_555,
output reg signed [15:0] RESULT_556,
output reg signed [15:0] RESULT_557,
output reg signed [15:0] RESULT_558,
output reg signed [15:0] RESULT_559,
output reg signed [15:0] RESULT_560,
output reg signed [15:0] RESULT_561,
output reg signed [15:0] RESULT_562,
output reg signed [15:0] RESULT_563,
output reg signed [15:0] RESULT_564,
output reg signed [15:0] RESULT_565,
output reg signed [15:0] RESULT_566,
output reg signed [15:0] RESULT_567,
output reg signed [15:0] RESULT_568,
output reg signed [15:0] RESULT_569,
output reg signed [15:0] RESULT_570,
output reg signed [15:0] RESULT_571,
output reg signed [15:0] RESULT_572,
output reg signed [15:0] RESULT_573,
output reg signed [15:0] RESULT_574,
output reg signed [15:0] RESULT_575,
output reg signed [15:0] RESULT_576,
output reg signed [15:0] RESULT_577,
output reg signed [15:0] RESULT_578,
output reg signed [15:0] RESULT_579,
output reg signed [15:0] RESULT_580,
output reg signed [15:0] RESULT_581,
output reg signed [15:0] RESULT_582,
output reg signed [15:0] RESULT_583,
output reg signed [15:0] RESULT_584,
output reg signed [15:0] RESULT_585,
output reg signed [15:0] RESULT_586,
output reg signed [15:0] RESULT_587,
output reg signed [15:0] RESULT_588,
output reg signed [15:0] RESULT_589,
output reg signed [15:0] RESULT_590,
output reg signed [15:0] RESULT_591,
output reg signed [15:0] RESULT_592,
output reg signed [15:0] RESULT_593,
output reg signed [15:0] RESULT_594,
output reg signed [15:0] RESULT_595,
output reg signed [15:0] RESULT_596,
output reg signed [15:0] RESULT_597,
output reg signed [15:0] RESULT_598,
output reg signed [15:0] RESULT_599,
output reg signed [15:0] RESULT_600,
output reg signed [15:0] RESULT_601,
output reg signed [15:0] RESULT_602,
output reg signed [15:0] RESULT_603,
output reg signed [15:0] RESULT_604,
output reg signed [15:0] RESULT_605,
output reg signed [15:0] RESULT_606,
output reg signed [15:0] RESULT_607,
output reg signed [15:0] RESULT_608,
output reg signed [15:0] RESULT_609,
output reg signed [15:0] RESULT_610,
output reg signed [15:0] RESULT_611,
output reg signed [15:0] RESULT_612,
output reg signed [15:0] RESULT_613,
output reg signed [15:0] RESULT_614,
output reg signed [15:0] RESULT_615,
output reg signed [15:0] RESULT_616,
output reg signed [15:0] RESULT_617,
output reg signed [15:0] RESULT_618,
output reg signed [15:0] RESULT_619,
output reg signed [15:0] RESULT_620,
output reg signed [15:0] RESULT_621,
output reg signed [15:0] RESULT_622,
output reg signed [15:0] RESULT_623,
output reg signed [15:0] RESULT_624,
output reg signed [15:0] RESULT_625,
output reg signed [15:0] RESULT_626,
output reg signed [15:0] RESULT_627,
output reg signed [15:0] RESULT_628,
output reg signed [15:0] RESULT_629,
output reg signed [15:0] RESULT_630,
output reg signed [15:0] RESULT_631,
output reg signed [15:0] RESULT_632,
output reg signed [15:0] RESULT_633,
output reg signed [15:0] RESULT_634,
output reg signed [15:0] RESULT_635,
output reg signed [15:0] RESULT_636,
output reg signed [15:0] RESULT_637,
output reg signed [15:0] RESULT_638,
output reg signed [15:0] RESULT_639,
output reg signed [15:0] RESULT_640,
output reg signed [15:0] RESULT_641,
output reg signed [15:0] RESULT_642,
output reg signed [15:0] RESULT_643,
output reg signed [15:0] RESULT_644,
output reg signed [15:0] RESULT_645,
output reg signed [15:0] RESULT_646,
output reg signed [15:0] RESULT_647,
output reg signed [15:0] RESULT_648,
output reg signed [15:0] RESULT_649,
output reg signed [15:0] RESULT_650,
output reg signed [15:0] RESULT_651,
output reg signed [15:0] RESULT_652,
output reg signed [15:0] RESULT_653,
output reg signed [15:0] RESULT_654,
output reg signed [15:0] RESULT_655,
output reg signed [15:0] RESULT_656,
output reg signed [15:0] RESULT_657,
output reg signed [15:0] RESULT_658,
output reg signed [15:0] RESULT_659,
output reg signed [15:0] RESULT_660,
output reg signed [15:0] RESULT_661,
output reg signed [15:0] RESULT_662,
output reg signed [15:0] RESULT_663,
output reg signed [15:0] RESULT_664,
output reg signed [15:0] RESULT_665,
output reg signed [15:0] RESULT_666,
output reg signed [15:0] RESULT_667,
output reg signed [15:0] RESULT_668,
output reg signed [15:0] RESULT_669,
output reg signed [15:0] RESULT_670,
output reg signed [15:0] RESULT_671,
output reg signed [15:0] RESULT_672,
output reg signed [15:0] RESULT_673,
output reg signed [15:0] RESULT_674,
output reg signed [15:0] RESULT_675,
output reg signed [15:0] RESULT_676,
output reg signed [15:0] RESULT_677,
output reg signed [15:0] RESULT_678,
output reg signed [15:0] RESULT_679,
output reg signed [15:0] RESULT_680,
output reg signed [15:0] RESULT_681,
output reg signed [15:0] RESULT_682,
output reg signed [15:0] RESULT_683,
output reg signed [15:0] RESULT_684,
output reg signed [15:0] RESULT_685,
output reg signed [15:0] RESULT_686,
output reg signed [15:0] RESULT_687,
output reg signed [15:0] RESULT_688,
output reg signed [15:0] RESULT_689,
output reg signed [15:0] RESULT_690,
output reg signed [15:0] RESULT_691,
output reg signed [15:0] RESULT_692,
output reg signed [15:0] RESULT_693,
output reg signed [15:0] RESULT_694,
output reg signed [15:0] RESULT_695,
output reg signed [15:0] RESULT_696,
output reg signed [15:0] RESULT_697,
output reg signed [15:0] RESULT_698,
output reg signed [15:0] RESULT_699,
output reg signed [15:0] RESULT_700,
output reg signed [15:0] RESULT_701,
output reg signed [15:0] RESULT_702,
output reg signed [15:0] RESULT_703,
output reg signed [15:0] RESULT_704,
output reg signed [15:0] RESULT_705,
output reg signed [15:0] RESULT_706,
output reg signed [15:0] RESULT_707,
output reg signed [15:0] RESULT_708,
output reg signed [15:0] RESULT_709,
output reg signed [15:0] RESULT_710,
output reg signed [15:0] RESULT_711,
output reg signed [15:0] RESULT_712,
output reg signed [15:0] RESULT_713,
output reg signed [15:0] RESULT_714,
output reg signed [15:0] RESULT_715,
output reg signed [15:0] RESULT_716,
output reg signed [15:0] RESULT_717,
output reg signed [15:0] RESULT_718,
output reg signed [15:0] RESULT_719,
output reg signed [15:0] RESULT_720,
output reg signed [15:0] RESULT_721,
output reg signed [15:0] RESULT_722,
output reg signed [15:0] RESULT_723,
output reg signed [15:0] RESULT_724,
output reg signed [15:0] RESULT_725,
output reg signed [15:0] RESULT_726,
output reg signed [15:0] RESULT_727,
output reg signed [15:0] RESULT_728,
output reg signed [15:0] RESULT_729,
output reg signed [15:0] RESULT_730,
output reg signed [15:0] RESULT_731,
output reg signed [15:0] RESULT_732,
output reg signed [15:0] RESULT_733,
output reg signed [15:0] RESULT_734,
output reg signed [15:0] RESULT_735,
output reg signed [15:0] RESULT_736,
output reg signed [15:0] RESULT_737,
output reg signed [15:0] RESULT_738,
output reg signed [15:0] RESULT_739,
output reg signed [15:0] RESULT_740,
output reg signed [15:0] RESULT_741,
output reg signed [15:0] RESULT_742,
output reg signed [15:0] RESULT_743,
output reg signed [15:0] RESULT_744,
output reg signed [15:0] RESULT_745,
output reg signed [15:0] RESULT_746,
output reg signed [15:0] RESULT_747,
output reg signed [15:0] RESULT_748,
output reg signed [15:0] RESULT_749,
output reg signed [15:0] RESULT_750,
output reg signed [15:0] RESULT_751,
output reg signed [15:0] RESULT_752,
output reg signed [15:0] RESULT_753,
output reg signed [15:0] RESULT_754,
output reg signed [15:0] RESULT_755,
output reg signed [15:0] RESULT_756,
output reg signed [15:0] RESULT_757,
output reg signed [15:0] RESULT_758,
output reg signed [15:0] RESULT_759,
output reg signed [15:0] RESULT_760,
output reg signed [15:0] RESULT_761,
output reg signed [15:0] RESULT_762,
output reg signed [15:0] RESULT_763,
output reg signed [15:0] RESULT_764,
output reg signed [15:0] RESULT_765,
output reg signed [15:0] RESULT_766,
output reg signed [15:0] RESULT_767,
output reg signed [15:0] RESULT_768,
output reg signed [15:0] RESULT_769,
output reg signed [15:0] RESULT_770,
output reg signed [15:0] RESULT_771,
output reg signed [15:0] RESULT_772,
output reg signed [15:0] RESULT_773,
output reg signed [15:0] RESULT_774,
output reg signed [15:0] RESULT_775,
output reg signed [15:0] RESULT_776,
output reg signed [15:0] RESULT_777,
output reg signed [15:0] RESULT_778,
output reg signed [15:0] RESULT_779,
output reg signed [15:0] RESULT_780,
output reg signed [15:0] RESULT_781,
output reg signed [15:0] RESULT_782,
output reg signed [15:0] RESULT_783,
output reg signed [15:0] RESULT_784,
output reg signed [15:0] RESULT_785,
output reg signed [15:0] RESULT_786,
output reg signed [15:0] RESULT_787,
output reg signed [15:0] RESULT_788,
output reg signed [15:0] RESULT_789,
output reg signed [15:0] RESULT_790,
output reg signed [15:0] RESULT_791,
output reg signed [15:0] RESULT_792,
output reg signed [15:0] RESULT_793,
output reg signed [15:0] RESULT_794,
output reg signed [15:0] RESULT_795,
output reg signed [15:0] RESULT_796,
output reg signed [15:0] RESULT_797,
output reg signed [15:0] RESULT_798,
output reg signed [15:0] RESULT_799,
output reg signed [15:0] RESULT_800,
output reg signed [15:0] RESULT_801,
output reg signed [15:0] RESULT_802,
output reg signed [15:0] RESULT_803,
output reg signed [15:0] RESULT_804,
output reg signed [15:0] RESULT_805,
output reg signed [15:0] RESULT_806,
output reg signed [15:0] RESULT_807,
output reg signed [15:0] RESULT_808,
output reg signed [15:0] RESULT_809,
output reg signed [15:0] RESULT_810,
output reg signed [15:0] RESULT_811,
output reg signed [15:0] RESULT_812,
output reg signed [15:0] RESULT_813,
output reg signed [15:0] RESULT_814,
output reg signed [15:0] RESULT_815,
output reg signed [15:0] RESULT_816,
output reg signed [15:0] RESULT_817,
output reg signed [15:0] RESULT_818,
output reg signed [15:0] RESULT_819,
output reg signed [15:0] RESULT_820,
output reg signed [15:0] RESULT_821,
output reg signed [15:0] RESULT_822,
output reg signed [15:0] RESULT_823,
output reg signed [15:0] RESULT_824,
output reg signed [15:0] RESULT_825,
output reg signed [15:0] RESULT_826,
output reg signed [15:0] RESULT_827,
output reg signed [15:0] RESULT_828,
output reg signed [15:0] RESULT_829,
output reg signed [15:0] RESULT_830,
output reg signed [15:0] RESULT_831,
output reg signed [15:0] RESULT_832,
output reg signed [15:0] RESULT_833,
output reg signed [15:0] RESULT_834,
output reg signed [15:0] RESULT_835,
output reg signed [15:0] RESULT_836,
output reg signed [15:0] RESULT_837,
output reg signed [15:0] RESULT_838,
output reg signed [15:0] RESULT_839,
output reg signed [15:0] RESULT_840,
output reg signed [15:0] RESULT_841,
output reg signed [15:0] RESULT_842,
output reg signed [15:0] RESULT_843,
output reg signed [15:0] RESULT_844,
output reg signed [15:0] RESULT_845,
output reg signed [15:0] RESULT_846,
output reg signed [15:0] RESULT_847,
output reg signed [15:0] RESULT_848,
output reg signed [15:0] RESULT_849,
output reg signed [15:0] RESULT_850,
output reg signed [15:0] RESULT_851,
output reg signed [15:0] RESULT_852,
output reg signed [15:0] RESULT_853,
output reg signed [15:0] RESULT_854,
output reg signed [15:0] RESULT_855,
output reg signed [15:0] RESULT_856,
output reg signed [15:0] RESULT_857,
output reg signed [15:0] RESULT_858,
output reg signed [15:0] RESULT_859,
output reg signed [15:0] RESULT_860,
output reg signed [15:0] RESULT_861,
output reg signed [15:0] RESULT_862,
output reg signed [15:0] RESULT_863,
output reg signed [15:0] RESULT_864,
output reg signed [15:0] RESULT_865,
output reg signed [15:0] RESULT_866,
output reg signed [15:0] RESULT_867,
output reg signed [15:0] RESULT_868,
output reg signed [15:0] RESULT_869,
output reg signed [15:0] RESULT_870,
output reg signed [15:0] RESULT_871,
output reg signed [15:0] RESULT_872,
output reg signed [15:0] RESULT_873,
output reg signed [15:0] RESULT_874,
output reg signed [15:0] RESULT_875,
output reg signed [15:0] RESULT_876,
output reg signed [15:0] RESULT_877,
output reg signed [15:0] RESULT_878,
output reg signed [15:0] RESULT_879,
output reg signed [15:0] RESULT_880,
output reg signed [15:0] RESULT_881,
output reg signed [15:0] RESULT_882,
output reg signed [15:0] RESULT_883,
output reg signed [15:0] RESULT_884,
output reg signed [15:0] RESULT_885,
output reg signed [15:0] RESULT_886,
output reg signed [15:0] RESULT_887,
output reg signed [15:0] RESULT_888,
output reg signed [15:0] RESULT_889,
output reg signed [15:0] RESULT_890,
output reg signed [15:0] RESULT_891,
output reg signed [15:0] RESULT_892,
output reg signed [15:0] RESULT_893,
output reg signed [15:0] RESULT_894,
output reg signed [15:0] RESULT_895

);

   reg [5:0] count;
   reg case_enable;

   always @(posedge CLK or negedge RSTN) begin
      if (!RSTN) begin
         RESULT_0 <= 16'b0;
         RESULT_1 <= 16'b0;
         RESULT_2 <= 16'b0;
         RESULT_3 <= 16'b0;
         RESULT_4 <= 16'b0;
         RESULT_5 <= 16'b0;
         RESULT_6 <= 16'b0;
         RESULT_7 <= 16'b0;
         RESULT_8 <= 16'b0;
         RESULT_9 <= 16'b0;
         RESULT_10 <= 16'b0;
         RESULT_11 <= 16'b0;
         RESULT_12 <= 16'b0;
         RESULT_13 <= 16'b0;
         RESULT_14 <= 16'b0;
         RESULT_15 <= 16'b0;
         RESULT_16 <= 16'b0;
         RESULT_17 <= 16'b0;
         RESULT_18 <= 16'b0;
         RESULT_19 <= 16'b0;
         RESULT_20 <= 16'b0;
         RESULT_21 <= 16'b0;
         RESULT_22 <= 16'b0;
         RESULT_23 <= 16'b0;
         RESULT_24 <= 16'b0;
         RESULT_25 <= 16'b0;
         RESULT_26 <= 16'b0;
         RESULT_27 <= 16'b0;
         RESULT_28 <= 16'b0;
         RESULT_29 <= 16'b0;
         RESULT_30 <= 16'b0;
         RESULT_31 <= 16'b0;
         RESULT_32 <= 16'b0;
         RESULT_33 <= 16'b0;
         RESULT_34 <= 16'b0;
         RESULT_35 <= 16'b0;
         RESULT_36 <= 16'b0;
         RESULT_37 <= 16'b0;
         RESULT_38 <= 16'b0;
         RESULT_39 <= 16'b0;
         RESULT_40 <= 16'b0;
         RESULT_41 <= 16'b0;
         RESULT_42 <= 16'b0;
         RESULT_43 <= 16'b0;
         RESULT_44 <= 16'b0;
         RESULT_45 <= 16'b0;
         RESULT_46 <= 16'b0;
         RESULT_47 <= 16'b0;
         RESULT_48 <= 16'b0;
         RESULT_49 <= 16'b0;
         RESULT_50 <= 16'b0;
         RESULT_51 <= 16'b0;
         RESULT_52 <= 16'b0;
         RESULT_53 <= 16'b0;
         RESULT_54 <= 16'b0;
         RESULT_55 <= 16'b0;
         RESULT_56 <= 16'b0;
         RESULT_57 <= 16'b0;
         RESULT_58 <= 16'b0;
         RESULT_59 <= 16'b0;
         RESULT_60 <= 16'b0;
         RESULT_61 <= 16'b0;
         RESULT_62 <= 16'b0;
         RESULT_63 <= 16'b0;
         RESULT_64 <= 16'b0;
         RESULT_65 <= 16'b0;
         RESULT_66 <= 16'b0;
         RESULT_67 <= 16'b0;
         RESULT_68 <= 16'b0;
         RESULT_69 <= 16'b0;
         RESULT_70 <= 16'b0;
         RESULT_71 <= 16'b0;
         RESULT_72 <= 16'b0;
         RESULT_73 <= 16'b0;
         RESULT_74 <= 16'b0;
         RESULT_75 <= 16'b0;
         RESULT_76 <= 16'b0;
         RESULT_77 <= 16'b0;
         RESULT_78 <= 16'b0;
         RESULT_79 <= 16'b0;
         RESULT_80 <= 16'b0;
         RESULT_81 <= 16'b0;
         RESULT_82 <= 16'b0;
         RESULT_83 <= 16'b0;
         RESULT_84 <= 16'b0;
         RESULT_85 <= 16'b0;
         RESULT_86 <= 16'b0;
         RESULT_87 <= 16'b0;
         RESULT_88 <= 16'b0;
         RESULT_89 <= 16'b0;
         RESULT_90 <= 16'b0;
         RESULT_91 <= 16'b0;
         RESULT_92 <= 16'b0;
         RESULT_93 <= 16'b0;
         RESULT_94 <= 16'b0;
         RESULT_95 <= 16'b0;
         RESULT_96 <= 16'b0;
         RESULT_97 <= 16'b0;
         RESULT_98 <= 16'b0;
         RESULT_99 <= 16'b0;
         RESULT_100 <= 16'b0;
         RESULT_101 <= 16'b0;
         RESULT_102 <= 16'b0;
         RESULT_103 <= 16'b0;
         RESULT_104 <= 16'b0;
         RESULT_105 <= 16'b0;
         RESULT_106 <= 16'b0;
         RESULT_107 <= 16'b0;
         RESULT_108 <= 16'b0;
         RESULT_109 <= 16'b0;
         RESULT_110 <= 16'b0;
         RESULT_111 <= 16'b0;
         RESULT_112 <= 16'b0;
         RESULT_113 <= 16'b0;
         RESULT_114 <= 16'b0;
         RESULT_115 <= 16'b0;
         RESULT_116 <= 16'b0;
         RESULT_117 <= 16'b0;
         RESULT_118 <= 16'b0;
         RESULT_119 <= 16'b0;
         RESULT_120 <= 16'b0;
         RESULT_121 <= 16'b0;
         RESULT_122 <= 16'b0;
         RESULT_123 <= 16'b0;
         RESULT_124 <= 16'b0;
         RESULT_125 <= 16'b0;
         RESULT_126 <= 16'b0;
         RESULT_127 <= 16'b0;
         RESULT_128 <= 16'b0;
         RESULT_129 <= 16'b0;
         RESULT_130 <= 16'b0;
         RESULT_131 <= 16'b0;
         RESULT_132 <= 16'b0;
         RESULT_133 <= 16'b0;
         RESULT_134 <= 16'b0;
         RESULT_135 <= 16'b0;
         RESULT_136 <= 16'b0;
         RESULT_137 <= 16'b0;
         RESULT_138 <= 16'b0;
         RESULT_139 <= 16'b0;
         RESULT_140 <= 16'b0;
         RESULT_141 <= 16'b0;
         RESULT_142 <= 16'b0;
         RESULT_143 <= 16'b0;
         RESULT_144 <= 16'b0;
         RESULT_145 <= 16'b0;
         RESULT_146 <= 16'b0;
         RESULT_147 <= 16'b0;
         RESULT_148 <= 16'b0;
         RESULT_149 <= 16'b0;
         RESULT_150 <= 16'b0;
         RESULT_151 <= 16'b0;
         RESULT_152 <= 16'b0;
         RESULT_153 <= 16'b0;
         RESULT_154 <= 16'b0;
         RESULT_155 <= 16'b0;
         RESULT_156 <= 16'b0;
         RESULT_157 <= 16'b0;
         RESULT_158 <= 16'b0;
         RESULT_159 <= 16'b0;
         RESULT_160 <= 16'b0;
         RESULT_161 <= 16'b0;
         RESULT_162 <= 16'b0;
         RESULT_163 <= 16'b0;
         RESULT_164 <= 16'b0;
         RESULT_165 <= 16'b0;
         RESULT_166 <= 16'b0;
         RESULT_167 <= 16'b0;
         RESULT_168 <= 16'b0;
         RESULT_169 <= 16'b0;
         RESULT_170 <= 16'b0;
         RESULT_171 <= 16'b0;
         RESULT_172 <= 16'b0;
         RESULT_173 <= 16'b0;
         RESULT_174 <= 16'b0;
         RESULT_175 <= 16'b0;
         RESULT_176 <= 16'b0;
         RESULT_177 <= 16'b0;
         RESULT_178 <= 16'b0;
         RESULT_179 <= 16'b0;
         RESULT_180 <= 16'b0;
         RESULT_181 <= 16'b0;
         RESULT_182 <= 16'b0;
         RESULT_183 <= 16'b0;
         RESULT_184 <= 16'b0;
         RESULT_185 <= 16'b0;
         RESULT_186 <= 16'b0;
         RESULT_187 <= 16'b0;
         RESULT_188 <= 16'b0;
         RESULT_189 <= 16'b0;
         RESULT_190 <= 16'b0;
         RESULT_191 <= 16'b0;
         RESULT_192 <= 16'b0;
         RESULT_193 <= 16'b0;
         RESULT_194 <= 16'b0;
         RESULT_195 <= 16'b0;
         RESULT_196 <= 16'b0;
         RESULT_197 <= 16'b0;
         RESULT_198 <= 16'b0;
         RESULT_199 <= 16'b0;
         RESULT_200 <= 16'b0;
         RESULT_201 <= 16'b0;
         RESULT_202 <= 16'b0;
         RESULT_203 <= 16'b0;
         RESULT_204 <= 16'b0;
         RESULT_205 <= 16'b0;
         RESULT_206 <= 16'b0;
         RESULT_207 <= 16'b0;
         RESULT_208 <= 16'b0;
         RESULT_209 <= 16'b0;
         RESULT_210 <= 16'b0;
         RESULT_211 <= 16'b0;
         RESULT_212 <= 16'b0;
         RESULT_213 <= 16'b0;
         RESULT_214 <= 16'b0;
         RESULT_215 <= 16'b0;
         RESULT_216 <= 16'b0;
         RESULT_217 <= 16'b0;
         RESULT_218 <= 16'b0;
         RESULT_219 <= 16'b0;
         RESULT_220 <= 16'b0;
         RESULT_221 <= 16'b0;
         RESULT_222 <= 16'b0;
         RESULT_223 <= 16'b0;
         RESULT_224 <= 16'b0;
         RESULT_225 <= 16'b0;
         RESULT_226 <= 16'b0;
         RESULT_227 <= 16'b0;
         RESULT_228 <= 16'b0;
         RESULT_229 <= 16'b0;
         RESULT_230 <= 16'b0;
         RESULT_231 <= 16'b0;
         RESULT_232 <= 16'b0;
         RESULT_233 <= 16'b0;
         RESULT_234 <= 16'b0;
         RESULT_235 <= 16'b0;
         RESULT_236 <= 16'b0;
         RESULT_237 <= 16'b0;
         RESULT_238 <= 16'b0;
         RESULT_239 <= 16'b0;
         RESULT_240 <= 16'b0;
         RESULT_241 <= 16'b0;
         RESULT_242 <= 16'b0;
         RESULT_243 <= 16'b0;
         RESULT_244 <= 16'b0;
         RESULT_245 <= 16'b0;
         RESULT_246 <= 16'b0;
         RESULT_247 <= 16'b0;
         RESULT_248 <= 16'b0;
         RESULT_249 <= 16'b0;
         RESULT_250 <= 16'b0;
         RESULT_251 <= 16'b0;
         RESULT_252 <= 16'b0;
         RESULT_253 <= 16'b0;
         RESULT_254 <= 16'b0;
         RESULT_255 <= 16'b0;
         RESULT_256 <= 16'b0;
         RESULT_257 <= 16'b0;
         RESULT_258 <= 16'b0;
         RESULT_259 <= 16'b0;
         RESULT_260 <= 16'b0;
         RESULT_261 <= 16'b0;
         RESULT_262 <= 16'b0;
         RESULT_263 <= 16'b0;
         RESULT_264 <= 16'b0;
         RESULT_265 <= 16'b0;
         RESULT_266 <= 16'b0;
         RESULT_267 <= 16'b0;
         RESULT_268 <= 16'b0;
         RESULT_269 <= 16'b0;
         RESULT_270 <= 16'b0;
         RESULT_271 <= 16'b0;
         RESULT_272 <= 16'b0;
         RESULT_273 <= 16'b0;
         RESULT_274 <= 16'b0;
         RESULT_275 <= 16'b0;
         RESULT_276 <= 16'b0;
         RESULT_277 <= 16'b0;
         RESULT_278 <= 16'b0;
         RESULT_279 <= 16'b0;
         RESULT_280 <= 16'b0;
         RESULT_281 <= 16'b0;
         RESULT_282 <= 16'b0;
         RESULT_283 <= 16'b0;
         RESULT_284 <= 16'b0;
         RESULT_285 <= 16'b0;
         RESULT_286 <= 16'b0;
         RESULT_287 <= 16'b0;
         RESULT_288 <= 16'b0;
         RESULT_289 <= 16'b0;
         RESULT_290 <= 16'b0;
         RESULT_291 <= 16'b0;
         RESULT_292 <= 16'b0;
         RESULT_293 <= 16'b0;
         RESULT_294 <= 16'b0;
         RESULT_295 <= 16'b0;
         RESULT_296 <= 16'b0;
         RESULT_297 <= 16'b0;
         RESULT_298 <= 16'b0;
         RESULT_299 <= 16'b0;
         RESULT_300 <= 16'b0;
         RESULT_301 <= 16'b0;
         RESULT_302 <= 16'b0;
         RESULT_303 <= 16'b0;
         RESULT_304 <= 16'b0;
         RESULT_305 <= 16'b0;
         RESULT_306 <= 16'b0;
         RESULT_307 <= 16'b0;
         RESULT_308 <= 16'b0;
         RESULT_309 <= 16'b0;
         RESULT_310 <= 16'b0;
         RESULT_311 <= 16'b0;
         RESULT_312 <= 16'b0;
         RESULT_313 <= 16'b0;
         RESULT_314 <= 16'b0;
         RESULT_315 <= 16'b0;
         RESULT_316 <= 16'b0;
         RESULT_317 <= 16'b0;
         RESULT_318 <= 16'b0;
         RESULT_319 <= 16'b0;
         RESULT_320 <= 16'b0;
         RESULT_321 <= 16'b0;
         RESULT_322 <= 16'b0;
         RESULT_323 <= 16'b0;
         RESULT_324 <= 16'b0;
         RESULT_325 <= 16'b0;
         RESULT_326 <= 16'b0;
         RESULT_327 <= 16'b0;
         RESULT_328 <= 16'b0;
         RESULT_329 <= 16'b0;
         RESULT_330 <= 16'b0;
         RESULT_331 <= 16'b0;
         RESULT_332 <= 16'b0;
         RESULT_333 <= 16'b0;
         RESULT_334 <= 16'b0;
         RESULT_335 <= 16'b0;
         RESULT_336 <= 16'b0;
         RESULT_337 <= 16'b0;
         RESULT_338 <= 16'b0;
         RESULT_339 <= 16'b0;
         RESULT_340 <= 16'b0;
         RESULT_341 <= 16'b0;
         RESULT_342 <= 16'b0;
         RESULT_343 <= 16'b0;
         RESULT_344 <= 16'b0;
         RESULT_345 <= 16'b0;
         RESULT_346 <= 16'b0;
         RESULT_347 <= 16'b0;
         RESULT_348 <= 16'b0;
         RESULT_349 <= 16'b0;
         RESULT_350 <= 16'b0;
         RESULT_351 <= 16'b0;
         RESULT_352 <= 16'b0;
         RESULT_353 <= 16'b0;
         RESULT_354 <= 16'b0;
         RESULT_355 <= 16'b0;
         RESULT_356 <= 16'b0;
         RESULT_357 <= 16'b0;
         RESULT_358 <= 16'b0;
         RESULT_359 <= 16'b0;
         RESULT_360 <= 16'b0;
         RESULT_361 <= 16'b0;
         RESULT_362 <= 16'b0;
         RESULT_363 <= 16'b0;
         RESULT_364 <= 16'b0;
         RESULT_365 <= 16'b0;
         RESULT_366 <= 16'b0;
         RESULT_367 <= 16'b0;
         RESULT_368 <= 16'b0;
         RESULT_369 <= 16'b0;
         RESULT_370 <= 16'b0;
         RESULT_371 <= 16'b0;
         RESULT_372 <= 16'b0;
         RESULT_373 <= 16'b0;
         RESULT_374 <= 16'b0;
         RESULT_375 <= 16'b0;
         RESULT_376 <= 16'b0;
         RESULT_377 <= 16'b0;
         RESULT_378 <= 16'b0;
         RESULT_379 <= 16'b0;
         RESULT_380 <= 16'b0;
         RESULT_381 <= 16'b0;
         RESULT_382 <= 16'b0;
         RESULT_383 <= 16'b0;
         RESULT_384 <= 16'b0;
         RESULT_385 <= 16'b0;
         RESULT_386 <= 16'b0;
         RESULT_387 <= 16'b0;
         RESULT_388 <= 16'b0;
         RESULT_389 <= 16'b0;
         RESULT_390 <= 16'b0;
         RESULT_391 <= 16'b0;
         RESULT_392 <= 16'b0;
         RESULT_393 <= 16'b0;
         RESULT_394 <= 16'b0;
         RESULT_395 <= 16'b0;
         RESULT_396 <= 16'b0;
         RESULT_397 <= 16'b0;
         RESULT_398 <= 16'b0;
         RESULT_399 <= 16'b0;
         RESULT_400 <= 16'b0;
         RESULT_401 <= 16'b0;
         RESULT_402 <= 16'b0;
         RESULT_403 <= 16'b0;
         RESULT_404 <= 16'b0;
         RESULT_405 <= 16'b0;
         RESULT_406 <= 16'b0;
         RESULT_407 <= 16'b0;
         RESULT_408 <= 16'b0;
         RESULT_409 <= 16'b0;
         RESULT_410 <= 16'b0;
         RESULT_411 <= 16'b0;
         RESULT_412 <= 16'b0;
         RESULT_413 <= 16'b0;
         RESULT_414 <= 16'b0;
         RESULT_415 <= 16'b0;
         RESULT_416 <= 16'b0;
         RESULT_417 <= 16'b0;
         RESULT_418 <= 16'b0;
         RESULT_419 <= 16'b0;
         RESULT_420 <= 16'b0;
         RESULT_421 <= 16'b0;
         RESULT_422 <= 16'b0;
         RESULT_423 <= 16'b0;
         RESULT_424 <= 16'b0;
         RESULT_425 <= 16'b0;
         RESULT_426 <= 16'b0;
         RESULT_427 <= 16'b0;
         RESULT_428 <= 16'b0;
         RESULT_429 <= 16'b0;
         RESULT_430 <= 16'b0;
         RESULT_431 <= 16'b0;
         RESULT_432 <= 16'b0;
         RESULT_433 <= 16'b0;
         RESULT_434 <= 16'b0;
         RESULT_435 <= 16'b0;
         RESULT_436 <= 16'b0;
         RESULT_437 <= 16'b0;
         RESULT_438 <= 16'b0;
         RESULT_439 <= 16'b0;
         RESULT_440 <= 16'b0;
         RESULT_441 <= 16'b0;
         RESULT_442 <= 16'b0;
         RESULT_443 <= 16'b0;
         RESULT_444 <= 16'b0;
         RESULT_445 <= 16'b0;
         RESULT_446 <= 16'b0;
         RESULT_447 <= 16'b0;
         RESULT_448 <= 16'b0;
         RESULT_449 <= 16'b0;
         RESULT_450 <= 16'b0;
         RESULT_451 <= 16'b0;
         RESULT_452 <= 16'b0;
         RESULT_453 <= 16'b0;
         RESULT_454 <= 16'b0;
         RESULT_455 <= 16'b0;
         RESULT_456 <= 16'b0;
         RESULT_457 <= 16'b0;
         RESULT_458 <= 16'b0;
         RESULT_459 <= 16'b0;
         RESULT_460 <= 16'b0;
         RESULT_461 <= 16'b0;
         RESULT_462 <= 16'b0;
         RESULT_463 <= 16'b0;
         RESULT_464 <= 16'b0;
         RESULT_465 <= 16'b0;
         RESULT_466 <= 16'b0;
         RESULT_467 <= 16'b0;
         RESULT_468 <= 16'b0;
         RESULT_469 <= 16'b0;
         RESULT_470 <= 16'b0;
         RESULT_471 <= 16'b0;
         RESULT_472 <= 16'b0;
         RESULT_473 <= 16'b0;
         RESULT_474 <= 16'b0;
         RESULT_475 <= 16'b0;
         RESULT_476 <= 16'b0;
         RESULT_477 <= 16'b0;
         RESULT_478 <= 16'b0;
         RESULT_479 <= 16'b0;
         RESULT_480 <= 16'b0;
         RESULT_481 <= 16'b0;
         RESULT_482 <= 16'b0;
         RESULT_483 <= 16'b0;
         RESULT_484 <= 16'b0;
         RESULT_485 <= 16'b0;
         RESULT_486 <= 16'b0;
         RESULT_487 <= 16'b0;
         RESULT_488 <= 16'b0;
         RESULT_489 <= 16'b0;
         RESULT_490 <= 16'b0;
         RESULT_491 <= 16'b0;
         RESULT_492 <= 16'b0;
         RESULT_493 <= 16'b0;
         RESULT_494 <= 16'b0;
         RESULT_495 <= 16'b0;
         RESULT_496 <= 16'b0;
         RESULT_497 <= 16'b0;
         RESULT_498 <= 16'b0;
         RESULT_499 <= 16'b0;
         RESULT_500 <= 16'b0;
         RESULT_501 <= 16'b0;
         RESULT_502 <= 16'b0;
         RESULT_503 <= 16'b0;
         RESULT_504 <= 16'b0;
         RESULT_505 <= 16'b0;
         RESULT_506 <= 16'b0;
         RESULT_507 <= 16'b0;
         RESULT_508 <= 16'b0;
         RESULT_509 <= 16'b0;
         RESULT_510 <= 16'b0;
         RESULT_511 <= 16'b0;
         RESULT_512 <= 16'b0;
         RESULT_513 <= 16'b0;
         RESULT_514 <= 16'b0;
         RESULT_515 <= 16'b0;
         RESULT_516 <= 16'b0;
         RESULT_517 <= 16'b0;
         RESULT_518 <= 16'b0;
         RESULT_519 <= 16'b0;
         RESULT_520 <= 16'b0;
         RESULT_521 <= 16'b0;
         RESULT_522 <= 16'b0;
         RESULT_523 <= 16'b0;
         RESULT_524 <= 16'b0;
         RESULT_525 <= 16'b0;
         RESULT_526 <= 16'b0;
         RESULT_527 <= 16'b0;
         RESULT_528 <= 16'b0;
         RESULT_529 <= 16'b0;
         RESULT_530 <= 16'b0;
         RESULT_531 <= 16'b0;
         RESULT_532 <= 16'b0;
         RESULT_533 <= 16'b0;
         RESULT_534 <= 16'b0;
         RESULT_535 <= 16'b0;
         RESULT_536 <= 16'b0;
         RESULT_537 <= 16'b0;
         RESULT_538 <= 16'b0;
         RESULT_539 <= 16'b0;
         RESULT_540 <= 16'b0;
         RESULT_541 <= 16'b0;
         RESULT_542 <= 16'b0;
         RESULT_543 <= 16'b0;
         RESULT_544 <= 16'b0;
         RESULT_545 <= 16'b0;
         RESULT_546 <= 16'b0;
         RESULT_547 <= 16'b0;
         RESULT_548 <= 16'b0;
         RESULT_549 <= 16'b0;
         RESULT_550 <= 16'b0;
         RESULT_551 <= 16'b0;
         RESULT_552 <= 16'b0;
         RESULT_553 <= 16'b0;
         RESULT_554 <= 16'b0;
         RESULT_555 <= 16'b0;
         RESULT_556 <= 16'b0;
         RESULT_557 <= 16'b0;
         RESULT_558 <= 16'b0;
         RESULT_559 <= 16'b0;
         RESULT_560 <= 16'b0;
         RESULT_561 <= 16'b0;
         RESULT_562 <= 16'b0;
         RESULT_563 <= 16'b0;
         RESULT_564 <= 16'b0;
         RESULT_565 <= 16'b0;
         RESULT_566 <= 16'b0;
         RESULT_567 <= 16'b0;
         RESULT_568 <= 16'b0;
         RESULT_569 <= 16'b0;
         RESULT_570 <= 16'b0;
         RESULT_571 <= 16'b0;
         RESULT_572 <= 16'b0;
         RESULT_573 <= 16'b0;
         RESULT_574 <= 16'b0;
         RESULT_575 <= 16'b0;
         RESULT_576 <= 16'b0;
         RESULT_577 <= 16'b0;
         RESULT_578 <= 16'b0;
         RESULT_579 <= 16'b0;
         RESULT_580 <= 16'b0;
         RESULT_581 <= 16'b0;
         RESULT_582 <= 16'b0;
         RESULT_583 <= 16'b0;
         RESULT_584 <= 16'b0;
         RESULT_585 <= 16'b0;
         RESULT_586 <= 16'b0;
         RESULT_587 <= 16'b0;
         RESULT_588 <= 16'b0;
         RESULT_589 <= 16'b0;
         RESULT_590 <= 16'b0;
         RESULT_591 <= 16'b0;
         RESULT_592 <= 16'b0;
         RESULT_593 <= 16'b0;
         RESULT_594 <= 16'b0;
         RESULT_595 <= 16'b0;
         RESULT_596 <= 16'b0;
         RESULT_597 <= 16'b0;
         RESULT_598 <= 16'b0;
         RESULT_599 <= 16'b0;
         RESULT_600 <= 16'b0;
         RESULT_601 <= 16'b0;
         RESULT_602 <= 16'b0;
         RESULT_603 <= 16'b0;
         RESULT_604 <= 16'b0;
         RESULT_605 <= 16'b0;
         RESULT_606 <= 16'b0;
         RESULT_607 <= 16'b0;
         RESULT_608 <= 16'b0;
         RESULT_609 <= 16'b0;
         RESULT_610 <= 16'b0;
         RESULT_611 <= 16'b0;
         RESULT_612 <= 16'b0;
         RESULT_613 <= 16'b0;
         RESULT_614 <= 16'b0;
         RESULT_615 <= 16'b0;
         RESULT_616 <= 16'b0;
         RESULT_617 <= 16'b0;
         RESULT_618 <= 16'b0;
         RESULT_619 <= 16'b0;
         RESULT_620 <= 16'b0;
         RESULT_621 <= 16'b0;
         RESULT_622 <= 16'b0;
         RESULT_623 <= 16'b0;
         RESULT_624 <= 16'b0;
         RESULT_625 <= 16'b0;
         RESULT_626 <= 16'b0;
         RESULT_627 <= 16'b0;
         RESULT_628 <= 16'b0;
         RESULT_629 <= 16'b0;
         RESULT_630 <= 16'b0;
         RESULT_631 <= 16'b0;
         RESULT_632 <= 16'b0;
         RESULT_633 <= 16'b0;
         RESULT_634 <= 16'b0;
         RESULT_635 <= 16'b0;
         RESULT_636 <= 16'b0;
         RESULT_637 <= 16'b0;
         RESULT_638 <= 16'b0;
         RESULT_639 <= 16'b0;
         RESULT_640 <= 16'b0;
         RESULT_641 <= 16'b0;
         RESULT_642 <= 16'b0;
         RESULT_643 <= 16'b0;
         RESULT_644 <= 16'b0;
         RESULT_645 <= 16'b0;
         RESULT_646 <= 16'b0;
         RESULT_647 <= 16'b0;
         RESULT_648 <= 16'b0;
         RESULT_649 <= 16'b0;
         RESULT_650 <= 16'b0;
         RESULT_651 <= 16'b0;
         RESULT_652 <= 16'b0;
         RESULT_653 <= 16'b0;
         RESULT_654 <= 16'b0;
         RESULT_655 <= 16'b0;
         RESULT_656 <= 16'b0;
         RESULT_657 <= 16'b0;
         RESULT_658 <= 16'b0;
         RESULT_659 <= 16'b0;
         RESULT_660 <= 16'b0;
         RESULT_661 <= 16'b0;
         RESULT_662 <= 16'b0;
         RESULT_663 <= 16'b0;
         RESULT_664 <= 16'b0;
         RESULT_665 <= 16'b0;
         RESULT_666 <= 16'b0;
         RESULT_667 <= 16'b0;
         RESULT_668 <= 16'b0;
         RESULT_669 <= 16'b0;
         RESULT_670 <= 16'b0;
         RESULT_671 <= 16'b0;
         RESULT_672 <= 16'b0;
         RESULT_673 <= 16'b0;
         RESULT_674 <= 16'b0;
         RESULT_675 <= 16'b0;
         RESULT_676 <= 16'b0;
         RESULT_677 <= 16'b0;
         RESULT_678 <= 16'b0;
         RESULT_679 <= 16'b0;
         RESULT_680 <= 16'b0;
         RESULT_681 <= 16'b0;
         RESULT_682 <= 16'b0;
         RESULT_683 <= 16'b0;
         RESULT_684 <= 16'b0;
         RESULT_685 <= 16'b0;
         RESULT_686 <= 16'b0;
         RESULT_687 <= 16'b0;
         RESULT_688 <= 16'b0;
         RESULT_689 <= 16'b0;
         RESULT_690 <= 16'b0;
         RESULT_691 <= 16'b0;
         RESULT_692 <= 16'b0;
         RESULT_693 <= 16'b0;
         RESULT_694 <= 16'b0;
         RESULT_695 <= 16'b0;
         RESULT_696 <= 16'b0;
         RESULT_697 <= 16'b0;
         RESULT_698 <= 16'b0;
         RESULT_699 <= 16'b0;
         RESULT_700 <= 16'b0;
         RESULT_701 <= 16'b0;
         RESULT_702 <= 16'b0;
         RESULT_703 <= 16'b0;
         RESULT_704 <= 16'b0;
         RESULT_705 <= 16'b0;
         RESULT_706 <= 16'b0;
         RESULT_707 <= 16'b0;
         RESULT_708 <= 16'b0;
         RESULT_709 <= 16'b0;
         RESULT_710 <= 16'b0;
         RESULT_711 <= 16'b0;
         RESULT_712 <= 16'b0;
         RESULT_713 <= 16'b0;
         RESULT_714 <= 16'b0;
         RESULT_715 <= 16'b0;
         RESULT_716 <= 16'b0;
         RESULT_717 <= 16'b0;
         RESULT_718 <= 16'b0;
         RESULT_719 <= 16'b0;
         RESULT_720 <= 16'b0;
         RESULT_721 <= 16'b0;
         RESULT_722 <= 16'b0;
         RESULT_723 <= 16'b0;
         RESULT_724 <= 16'b0;
         RESULT_725 <= 16'b0;
         RESULT_726 <= 16'b0;
         RESULT_727 <= 16'b0;
         RESULT_728 <= 16'b0;
         RESULT_729 <= 16'b0;
         RESULT_730 <= 16'b0;
         RESULT_731 <= 16'b0;
         RESULT_732 <= 16'b0;
         RESULT_733 <= 16'b0;
         RESULT_734 <= 16'b0;
         RESULT_735 <= 16'b0;
         RESULT_736 <= 16'b0;
         RESULT_737 <= 16'b0;
         RESULT_738 <= 16'b0;
         RESULT_739 <= 16'b0;
         RESULT_740 <= 16'b0;
         RESULT_741 <= 16'b0;
         RESULT_742 <= 16'b0;
         RESULT_743 <= 16'b0;
         RESULT_744 <= 16'b0;
         RESULT_745 <= 16'b0;
         RESULT_746 <= 16'b0;
         RESULT_747 <= 16'b0;
         RESULT_748 <= 16'b0;
         RESULT_749 <= 16'b0;
         RESULT_750 <= 16'b0;
         RESULT_751 <= 16'b0;
         RESULT_752 <= 16'b0;
         RESULT_753 <= 16'b0;
         RESULT_754 <= 16'b0;
         RESULT_755 <= 16'b0;
         RESULT_756 <= 16'b0;
         RESULT_757 <= 16'b0;
         RESULT_758 <= 16'b0;
         RESULT_759 <= 16'b0;
         RESULT_760 <= 16'b0;
         RESULT_761 <= 16'b0;
         RESULT_762 <= 16'b0;
         RESULT_763 <= 16'b0;
         RESULT_764 <= 16'b0;
         RESULT_765 <= 16'b0;
         RESULT_766 <= 16'b0;
         RESULT_767 <= 16'b0;
         RESULT_768 <= 16'b0;
         RESULT_769 <= 16'b0;
         RESULT_770 <= 16'b0;
         RESULT_771 <= 16'b0;
         RESULT_772 <= 16'b0;
         RESULT_773 <= 16'b0;
         RESULT_774 <= 16'b0;
         RESULT_775 <= 16'b0;
         RESULT_776 <= 16'b0;
         RESULT_777 <= 16'b0;
         RESULT_778 <= 16'b0;
         RESULT_779 <= 16'b0;
         RESULT_780 <= 16'b0;
         RESULT_781 <= 16'b0;
         RESULT_782 <= 16'b0;
         RESULT_783 <= 16'b0;
         RESULT_784 <= 16'b0;
         RESULT_785 <= 16'b0;
         RESULT_786 <= 16'b0;
         RESULT_787 <= 16'b0;
         RESULT_788 <= 16'b0;
         RESULT_789 <= 16'b0;
         RESULT_790 <= 16'b0;
         RESULT_791 <= 16'b0;
         RESULT_792 <= 16'b0;
         RESULT_793 <= 16'b0;
         RESULT_794 <= 16'b0;
         RESULT_795 <= 16'b0;
         RESULT_796 <= 16'b0;
         RESULT_797 <= 16'b0;
         RESULT_798 <= 16'b0;
         RESULT_799 <= 16'b0;
         RESULT_800 <= 16'b0;
         RESULT_801 <= 16'b0;
         RESULT_802 <= 16'b0;
         RESULT_803 <= 16'b0;
         RESULT_804 <= 16'b0;
         RESULT_805 <= 16'b0;
         RESULT_806 <= 16'b0;
         RESULT_807 <= 16'b0;
         RESULT_808 <= 16'b0;
         RESULT_809 <= 16'b0;
         RESULT_810 <= 16'b0;
         RESULT_811 <= 16'b0;
         RESULT_812 <= 16'b0;
         RESULT_813 <= 16'b0;
         RESULT_814 <= 16'b0;
         RESULT_815 <= 16'b0;
         RESULT_816 <= 16'b0;
         RESULT_817 <= 16'b0;
         RESULT_818 <= 16'b0;
         RESULT_819 <= 16'b0;
         RESULT_820 <= 16'b0;
         RESULT_821 <= 16'b0;
         RESULT_822 <= 16'b0;
         RESULT_823 <= 16'b0;
         RESULT_824 <= 16'b0;
         RESULT_825 <= 16'b0;
         RESULT_826 <= 16'b0;
         RESULT_827 <= 16'b0;
         RESULT_828 <= 16'b0;
         RESULT_829 <= 16'b0;
         RESULT_830 <= 16'b0;
         RESULT_831 <= 16'b0;
         RESULT_832 <= 16'b0;
         RESULT_833 <= 16'b0;
         RESULT_834 <= 16'b0;
         RESULT_835 <= 16'b0;
         RESULT_836 <= 16'b0;
         RESULT_837 <= 16'b0;
         RESULT_838 <= 16'b0;
         RESULT_839 <= 16'b0;
         RESULT_840 <= 16'b0;
         RESULT_841 <= 16'b0;
         RESULT_842 <= 16'b0;
         RESULT_843 <= 16'b0;
         RESULT_844 <= 16'b0;
         RESULT_845 <= 16'b0;
         RESULT_846 <= 16'b0;
         RESULT_847 <= 16'b0;
         RESULT_848 <= 16'b0;
         RESULT_849 <= 16'b0;
         RESULT_850 <= 16'b0;
         RESULT_851 <= 16'b0;
         RESULT_852 <= 16'b0;
         RESULT_853 <= 16'b0;
         RESULT_854 <= 16'b0;
         RESULT_855 <= 16'b0;
         RESULT_856 <= 16'b0;
         RESULT_857 <= 16'b0;
         RESULT_858 <= 16'b0;
         RESULT_859 <= 16'b0;
         RESULT_860 <= 16'b0;
         RESULT_861 <= 16'b0;
         RESULT_862 <= 16'b0;
         RESULT_863 <= 16'b0;
         RESULT_864 <= 16'b0;
         RESULT_865 <= 16'b0;
         RESULT_866 <= 16'b0;
         RESULT_867 <= 16'b0;
         RESULT_868 <= 16'b0;
         RESULT_869 <= 16'b0;
         RESULT_870 <= 16'b0;
         RESULT_871 <= 16'b0;
         RESULT_872 <= 16'b0;
         RESULT_873 <= 16'b0;
         RESULT_874 <= 16'b0;
         RESULT_875 <= 16'b0;
         RESULT_876 <= 16'b0;
         RESULT_877 <= 16'b0;
         RESULT_878 <= 16'b0;
         RESULT_879 <= 16'b0;
         RESULT_880 <= 16'b0;
         RESULT_881 <= 16'b0;
         RESULT_882 <= 16'b0;
         RESULT_883 <= 16'b0;
         RESULT_884 <= 16'b0;
         RESULT_885 <= 16'b0;
         RESULT_886 <= 16'b0;
         RESULT_887 <= 16'b0;
         RESULT_888 <= 16'b0;
         RESULT_889 <= 16'b0;
         RESULT_890 <= 16'b0;
         RESULT_891 <= 16'b0;
         RESULT_892 <= 16'b0;
         RESULT_893 <= 16'b0;
         RESULT_894 <= 16'b0;
         RESULT_895 <= 16'b0;
      end else if(case_enable) begin
         case (count)
			3: begin
			RESULT_192 <= RESULT_P18;
			end
			4: begin
			RESULT_193 <= RESULT_P18;
			RESULT_160 <= RESULT_P17;
			RESULT_384 <= RESULT_P28;
			end
			5: begin
			RESULT_194 <= RESULT_P18;
			RESULT_161 <= RESULT_P17;
			RESULT_385 <= RESULT_P28;
			RESULT_128 <= RESULT_P16;
			RESULT_352 <= RESULT_P27;
			RESULT_544 <= RESULT_P38;
			end
			6: begin
			RESULT_195 <= RESULT_P18;
			RESULT_162 <= RESULT_P17;
			RESULT_386 <= RESULT_P28;
			RESULT_129 <= RESULT_P16;
			RESULT_353 <= RESULT_P27;
			RESULT_545 <= RESULT_P38;
			RESULT_96 <= RESULT_P15;
			RESULT_320 <= RESULT_P26;
			RESULT_512 <= RESULT_P37;
			RESULT_672 <= RESULT_P48;
			end
			7: begin
			RESULT_196 <= RESULT_P18;
			RESULT_163 <= RESULT_P17;
			RESULT_387 <= RESULT_P28;
			RESULT_130 <= RESULT_P16;
			RESULT_354 <= RESULT_P27;
			RESULT_546 <= RESULT_P38;
			RESULT_97 <= RESULT_P15;
			RESULT_321 <= RESULT_P26;
			RESULT_513 <= RESULT_P37;
			RESULT_673 <= RESULT_P48;
			RESULT_64 <= RESULT_P14;
			RESULT_288 <= RESULT_P25;
			RESULT_480 <= RESULT_P36;
			RESULT_640 <= RESULT_P47;
			RESULT_768 <= RESULT_P58;
			end
			8: begin
			RESULT_197 <= RESULT_P18;
			RESULT_164 <= RESULT_P17;
			RESULT_388 <= RESULT_P28;
			RESULT_131 <= RESULT_P16;
			RESULT_355 <= RESULT_P27;
			RESULT_547 <= RESULT_P38;
			RESULT_98 <= RESULT_P15;
			RESULT_322 <= RESULT_P26;
			RESULT_514 <= RESULT_P37;
			RESULT_674 <= RESULT_P48;
			RESULT_65 <= RESULT_P14;
			RESULT_289 <= RESULT_P25;
			RESULT_481 <= RESULT_P36;
			RESULT_641 <= RESULT_P47;
			RESULT_769 <= RESULT_P58;
			RESULT_32 <= RESULT_P13;
			RESULT_256 <= RESULT_P24;
			RESULT_448 <= RESULT_P35;
			RESULT_608 <= RESULT_P46;
			RESULT_736 <= RESULT_P57;
			RESULT_832 <= RESULT_P68;
			end
			9: begin
			RESULT_198 <= RESULT_P18;
			RESULT_165 <= RESULT_P17;
			RESULT_389 <= RESULT_P28;
			RESULT_132 <= RESULT_P16;
			RESULT_356 <= RESULT_P27;
			RESULT_548 <= RESULT_P38;
			RESULT_99 <= RESULT_P15;
			RESULT_323 <= RESULT_P26;
			RESULT_515 <= RESULT_P37;
			RESULT_675 <= RESULT_P48;
			RESULT_66 <= RESULT_P14;
			RESULT_290 <= RESULT_P25;
			RESULT_482 <= RESULT_P36;
			RESULT_642 <= RESULT_P47;
			RESULT_770 <= RESULT_P58;
			RESULT_33 <= RESULT_P13;
			RESULT_257 <= RESULT_P24;
			RESULT_449 <= RESULT_P35;
			RESULT_609 <= RESULT_P46;
			RESULT_737 <= RESULT_P57;
			RESULT_833 <= RESULT_P68;
			RESULT_0 <= RESULT_P12;
			RESULT_224 <= RESULT_P23;
			RESULT_416 <= RESULT_P34;
			RESULT_576 <= RESULT_P45;
			RESULT_704 <= RESULT_P56;
			RESULT_800 <= RESULT_P67;
			RESULT_864 <= RESULT_P78;
			end
			10: begin
			RESULT_199 <= RESULT_P18;
			RESULT_166 <= RESULT_P17;
			RESULT_390 <= RESULT_P28;
			RESULT_133 <= RESULT_P16;
			RESULT_357 <= RESULT_P27;
			RESULT_549 <= RESULT_P38;
			RESULT_100 <= RESULT_P15;
			RESULT_324 <= RESULT_P26;
			RESULT_516 <= RESULT_P37;
			RESULT_676 <= RESULT_P48;
			RESULT_67 <= RESULT_P14;
			RESULT_291 <= RESULT_P25;
			RESULT_483 <= RESULT_P36;
			RESULT_643 <= RESULT_P47;
			RESULT_771 <= RESULT_P58;
			RESULT_34 <= RESULT_P13;
			RESULT_258 <= RESULT_P24;
			RESULT_450 <= RESULT_P35;
			RESULT_610 <= RESULT_P46;
			RESULT_738 <= RESULT_P57;
			RESULT_834 <= RESULT_P68;
			RESULT_1 <= RESULT_P12;
			RESULT_225 <= RESULT_P23;
			RESULT_417 <= RESULT_P34;
			RESULT_577 <= RESULT_P45;
			RESULT_705 <= RESULT_P56;
			RESULT_801 <= RESULT_P67;
			RESULT_865 <= RESULT_P78;
			end
			11: begin
			RESULT_200 <= RESULT_P18;
			RESULT_167 <= RESULT_P17;
			RESULT_391 <= RESULT_P28;
			RESULT_134 <= RESULT_P16;
			RESULT_358 <= RESULT_P27;
			RESULT_550 <= RESULT_P38;
			RESULT_101 <= RESULT_P15;
			RESULT_325 <= RESULT_P26;
			RESULT_517 <= RESULT_P37;
			RESULT_677 <= RESULT_P48;
			RESULT_68 <= RESULT_P14;
			RESULT_292 <= RESULT_P25;
			RESULT_484 <= RESULT_P36;
			RESULT_644 <= RESULT_P47;
			RESULT_772 <= RESULT_P58;
			RESULT_35 <= RESULT_P13;
			RESULT_259 <= RESULT_P24;
			RESULT_451 <= RESULT_P35;
			RESULT_611 <= RESULT_P46;
			RESULT_739 <= RESULT_P57;
			RESULT_835 <= RESULT_P68;
			RESULT_2 <= RESULT_P12;
			RESULT_226 <= RESULT_P23;
			RESULT_418 <= RESULT_P34;
			RESULT_578 <= RESULT_P45;
			RESULT_706 <= RESULT_P56;
			RESULT_802 <= RESULT_P67;
			RESULT_866 <= RESULT_P78;
			end
			12: begin
			RESULT_201 <= RESULT_P18;
			RESULT_168 <= RESULT_P17;
			RESULT_392 <= RESULT_P28;
			RESULT_135 <= RESULT_P16;
			RESULT_359 <= RESULT_P27;
			RESULT_551 <= RESULT_P38;
			RESULT_102 <= RESULT_P15;
			RESULT_326 <= RESULT_P26;
			RESULT_518 <= RESULT_P37;
			RESULT_678 <= RESULT_P48;
			RESULT_69 <= RESULT_P14;
			RESULT_293 <= RESULT_P25;
			RESULT_485 <= RESULT_P36;
			RESULT_645 <= RESULT_P47;
			RESULT_773 <= RESULT_P58;
			RESULT_36 <= RESULT_P13;
			RESULT_260 <= RESULT_P24;
			RESULT_452 <= RESULT_P35;
			RESULT_612 <= RESULT_P46;
			RESULT_740 <= RESULT_P57;
			RESULT_836 <= RESULT_P68;
			RESULT_3 <= RESULT_P12;
			RESULT_227 <= RESULT_P23;
			RESULT_419 <= RESULT_P34;
			RESULT_579 <= RESULT_P45;
			RESULT_707 <= RESULT_P56;
			RESULT_803 <= RESULT_P67;
			RESULT_867 <= RESULT_P78;
			end
			13: begin
			RESULT_202 <= RESULT_P18;
			RESULT_169 <= RESULT_P17;
			RESULT_393 <= RESULT_P28;
			RESULT_136 <= RESULT_P16;
			RESULT_360 <= RESULT_P27;
			RESULT_552 <= RESULT_P38;
			RESULT_103 <= RESULT_P15;
			RESULT_327 <= RESULT_P26;
			RESULT_519 <= RESULT_P37;
			RESULT_679 <= RESULT_P48;
			RESULT_70 <= RESULT_P14;
			RESULT_294 <= RESULT_P25;
			RESULT_486 <= RESULT_P36;
			RESULT_646 <= RESULT_P47;
			RESULT_774 <= RESULT_P58;
			RESULT_37 <= RESULT_P13;
			RESULT_261 <= RESULT_P24;
			RESULT_453 <= RESULT_P35;
			RESULT_613 <= RESULT_P46;
			RESULT_741 <= RESULT_P57;
			RESULT_837 <= RESULT_P68;
			RESULT_4 <= RESULT_P12;
			RESULT_228 <= RESULT_P23;
			RESULT_420 <= RESULT_P34;
			RESULT_580 <= RESULT_P45;
			RESULT_708 <= RESULT_P56;
			RESULT_804 <= RESULT_P67;
			RESULT_868 <= RESULT_P78;
			end
			14: begin
			RESULT_203 <= RESULT_P18;
			RESULT_170 <= RESULT_P17;
			RESULT_394 <= RESULT_P28;
			RESULT_137 <= RESULT_P16;
			RESULT_361 <= RESULT_P27;
			RESULT_553 <= RESULT_P38;
			RESULT_104 <= RESULT_P15;
			RESULT_328 <= RESULT_P26;
			RESULT_520 <= RESULT_P37;
			RESULT_680 <= RESULT_P48;
			RESULT_71 <= RESULT_P14;
			RESULT_295 <= RESULT_P25;
			RESULT_487 <= RESULT_P36;
			RESULT_647 <= RESULT_P47;
			RESULT_775 <= RESULT_P58;
			RESULT_38 <= RESULT_P13;
			RESULT_262 <= RESULT_P24;
			RESULT_454 <= RESULT_P35;
			RESULT_614 <= RESULT_P46;
			RESULT_742 <= RESULT_P57;
			RESULT_838 <= RESULT_P68;
			RESULT_5 <= RESULT_P12;
			RESULT_229 <= RESULT_P23;
			RESULT_421 <= RESULT_P34;
			RESULT_581 <= RESULT_P45;
			RESULT_709 <= RESULT_P56;
			RESULT_805 <= RESULT_P67;
			RESULT_869 <= RESULT_P78;
			end
			15: begin
			RESULT_204 <= RESULT_P18;
			RESULT_171 <= RESULT_P17;
			RESULT_395 <= RESULT_P28;
			RESULT_138 <= RESULT_P16;
			RESULT_362 <= RESULT_P27;
			RESULT_554 <= RESULT_P38;
			RESULT_105 <= RESULT_P15;
			RESULT_329 <= RESULT_P26;
			RESULT_521 <= RESULT_P37;
			RESULT_681 <= RESULT_P48;
			RESULT_72 <= RESULT_P14;
			RESULT_296 <= RESULT_P25;
			RESULT_488 <= RESULT_P36;
			RESULT_648 <= RESULT_P47;
			RESULT_776 <= RESULT_P58;
			RESULT_39 <= RESULT_P13;
			RESULT_263 <= RESULT_P24;
			RESULT_455 <= RESULT_P35;
			RESULT_615 <= RESULT_P46;
			RESULT_743 <= RESULT_P57;
			RESULT_839 <= RESULT_P68;
			RESULT_6 <= RESULT_P12;
			RESULT_230 <= RESULT_P23;
			RESULT_422 <= RESULT_P34;
			RESULT_582 <= RESULT_P45;
			RESULT_710 <= RESULT_P56;
			RESULT_806 <= RESULT_P67;
			RESULT_870 <= RESULT_P78;
			end
			16: begin
			RESULT_205 <= RESULT_P18;
			RESULT_172 <= RESULT_P17;
			RESULT_396 <= RESULT_P28;
			RESULT_139 <= RESULT_P16;
			RESULT_363 <= RESULT_P27;
			RESULT_555 <= RESULT_P38;
			RESULT_106 <= RESULT_P15;
			RESULT_330 <= RESULT_P26;
			RESULT_522 <= RESULT_P37;
			RESULT_682 <= RESULT_P48;
			RESULT_73 <= RESULT_P14;
			RESULT_297 <= RESULT_P25;
			RESULT_489 <= RESULT_P36;
			RESULT_649 <= RESULT_P47;
			RESULT_777 <= RESULT_P58;
			RESULT_40 <= RESULT_P13;
			RESULT_264 <= RESULT_P24;
			RESULT_456 <= RESULT_P35;
			RESULT_616 <= RESULT_P46;
			RESULT_744 <= RESULT_P57;
			RESULT_840 <= RESULT_P68;
			RESULT_7 <= RESULT_P12;
			RESULT_231 <= RESULT_P23;
			RESULT_423 <= RESULT_P34;
			RESULT_583 <= RESULT_P45;
			RESULT_711 <= RESULT_P56;
			RESULT_807 <= RESULT_P67;
			RESULT_871 <= RESULT_P78;
			end
			17: begin
			RESULT_206 <= RESULT_P18;
			RESULT_173 <= RESULT_P17;
			RESULT_397 <= RESULT_P28;
			RESULT_140 <= RESULT_P16;
			RESULT_364 <= RESULT_P27;
			RESULT_556 <= RESULT_P38;
			RESULT_107 <= RESULT_P15;
			RESULT_331 <= RESULT_P26;
			RESULT_523 <= RESULT_P37;
			RESULT_683 <= RESULT_P48;
			RESULT_74 <= RESULT_P14;
			RESULT_298 <= RESULT_P25;
			RESULT_490 <= RESULT_P36;
			RESULT_650 <= RESULT_P47;
			RESULT_778 <= RESULT_P58;
			RESULT_41 <= RESULT_P13;
			RESULT_265 <= RESULT_P24;
			RESULT_457 <= RESULT_P35;
			RESULT_617 <= RESULT_P46;
			RESULT_745 <= RESULT_P57;
			RESULT_841 <= RESULT_P68;
			RESULT_8 <= RESULT_P12;
			RESULT_232 <= RESULT_P23;
			RESULT_424 <= RESULT_P34;
			RESULT_584 <= RESULT_P45;
			RESULT_712 <= RESULT_P56;
			RESULT_808 <= RESULT_P67;
			RESULT_872 <= RESULT_P78;
			end
			18: begin
			RESULT_207 <= RESULT_P18;
			RESULT_174 <= RESULT_P17;
			RESULT_398 <= RESULT_P28;
			RESULT_141 <= RESULT_P16;
			RESULT_365 <= RESULT_P27;
			RESULT_557 <= RESULT_P38;
			RESULT_108 <= RESULT_P15;
			RESULT_332 <= RESULT_P26;
			RESULT_524 <= RESULT_P37;
			RESULT_684 <= RESULT_P48;
			RESULT_75 <= RESULT_P14;
			RESULT_299 <= RESULT_P25;
			RESULT_491 <= RESULT_P36;
			RESULT_651 <= RESULT_P47;
			RESULT_779 <= RESULT_P58;
			RESULT_42 <= RESULT_P13;
			RESULT_266 <= RESULT_P24;
			RESULT_458 <= RESULT_P35;
			RESULT_618 <= RESULT_P46;
			RESULT_746 <= RESULT_P57;
			RESULT_842 <= RESULT_P68;
			RESULT_9 <= RESULT_P12;
			RESULT_233 <= RESULT_P23;
			RESULT_425 <= RESULT_P34;
			RESULT_585 <= RESULT_P45;
			RESULT_713 <= RESULT_P56;
			RESULT_809 <= RESULT_P67;
			RESULT_873 <= RESULT_P78;
			end
			19: begin
			RESULT_208 <= RESULT_P18;
			RESULT_175 <= RESULT_P17;
			RESULT_399 <= RESULT_P28;
			RESULT_142 <= RESULT_P16;
			RESULT_366 <= RESULT_P27;
			RESULT_558 <= RESULT_P38;
			RESULT_109 <= RESULT_P15;
			RESULT_333 <= RESULT_P26;
			RESULT_525 <= RESULT_P37;
			RESULT_685 <= RESULT_P48;
			RESULT_76 <= RESULT_P14;
			RESULT_300 <= RESULT_P25;
			RESULT_492 <= RESULT_P36;
			RESULT_652 <= RESULT_P47;
			RESULT_780 <= RESULT_P58;
			RESULT_43 <= RESULT_P13;
			RESULT_267 <= RESULT_P24;
			RESULT_459 <= RESULT_P35;
			RESULT_619 <= RESULT_P46;
			RESULT_747 <= RESULT_P57;
			RESULT_843 <= RESULT_P68;
			RESULT_10 <= RESULT_P12;
			RESULT_234 <= RESULT_P23;
			RESULT_426 <= RESULT_P34;
			RESULT_586 <= RESULT_P45;
			RESULT_714 <= RESULT_P56;
			RESULT_810 <= RESULT_P67;
			RESULT_874 <= RESULT_P78;
			end
			20: begin
			RESULT_209 <= RESULT_P18;
			RESULT_176 <= RESULT_P17;
			RESULT_400 <= RESULT_P28;
			RESULT_143 <= RESULT_P16;
			RESULT_367 <= RESULT_P27;
			RESULT_559 <= RESULT_P38;
			RESULT_110 <= RESULT_P15;
			RESULT_334 <= RESULT_P26;
			RESULT_526 <= RESULT_P37;
			RESULT_686 <= RESULT_P48;
			RESULT_77 <= RESULT_P14;
			RESULT_301 <= RESULT_P25;
			RESULT_493 <= RESULT_P36;
			RESULT_653 <= RESULT_P47;
			RESULT_781 <= RESULT_P58;
			RESULT_44 <= RESULT_P13;
			RESULT_268 <= RESULT_P24;
			RESULT_460 <= RESULT_P35;
			RESULT_620 <= RESULT_P46;
			RESULT_748 <= RESULT_P57;
			RESULT_844 <= RESULT_P68;
			RESULT_11 <= RESULT_P12;
			RESULT_235 <= RESULT_P23;
			RESULT_427 <= RESULT_P34;
			RESULT_587 <= RESULT_P45;
			RESULT_715 <= RESULT_P56;
			RESULT_811 <= RESULT_P67;
			RESULT_875 <= RESULT_P78;
			end
			21: begin
			RESULT_210 <= RESULT_P18;
			RESULT_177 <= RESULT_P17;
			RESULT_401 <= RESULT_P28;
			RESULT_144 <= RESULT_P16;
			RESULT_368 <= RESULT_P27;
			RESULT_560 <= RESULT_P38;
			RESULT_111 <= RESULT_P15;
			RESULT_335 <= RESULT_P26;
			RESULT_527 <= RESULT_P37;
			RESULT_687 <= RESULT_P48;
			RESULT_78 <= RESULT_P14;
			RESULT_302 <= RESULT_P25;
			RESULT_494 <= RESULT_P36;
			RESULT_654 <= RESULT_P47;
			RESULT_782 <= RESULT_P58;
			RESULT_45 <= RESULT_P13;
			RESULT_269 <= RESULT_P24;
			RESULT_461 <= RESULT_P35;
			RESULT_621 <= RESULT_P46;
			RESULT_749 <= RESULT_P57;
			RESULT_845 <= RESULT_P68;
			RESULT_12 <= RESULT_P12;
			RESULT_236 <= RESULT_P23;
			RESULT_428 <= RESULT_P34;
			RESULT_588 <= RESULT_P45;
			RESULT_716 <= RESULT_P56;
			RESULT_812 <= RESULT_P67;
			RESULT_876 <= RESULT_P78;
			end
			22: begin
			RESULT_211 <= RESULT_P18;
			RESULT_178 <= RESULT_P17;
			RESULT_402 <= RESULT_P28;
			RESULT_145 <= RESULT_P16;
			RESULT_369 <= RESULT_P27;
			RESULT_561 <= RESULT_P38;
			RESULT_112 <= RESULT_P15;
			RESULT_336 <= RESULT_P26;
			RESULT_528 <= RESULT_P37;
			RESULT_688 <= RESULT_P48;
			RESULT_79 <= RESULT_P14;
			RESULT_303 <= RESULT_P25;
			RESULT_495 <= RESULT_P36;
			RESULT_655 <= RESULT_P47;
			RESULT_783 <= RESULT_P58;
			RESULT_46 <= RESULT_P13;
			RESULT_270 <= RESULT_P24;
			RESULT_462 <= RESULT_P35;
			RESULT_622 <= RESULT_P46;
			RESULT_750 <= RESULT_P57;
			RESULT_846 <= RESULT_P68;
			RESULT_13 <= RESULT_P12;
			RESULT_237 <= RESULT_P23;
			RESULT_429 <= RESULT_P34;
			RESULT_589 <= RESULT_P45;
			RESULT_717 <= RESULT_P56;
			RESULT_813 <= RESULT_P67;
			RESULT_877 <= RESULT_P78;
			end
			23: begin
			RESULT_212 <= RESULT_P18;
			RESULT_179 <= RESULT_P17;
			RESULT_403 <= RESULT_P28;
			RESULT_146 <= RESULT_P16;
			RESULT_370 <= RESULT_P27;
			RESULT_562 <= RESULT_P38;
			RESULT_113 <= RESULT_P15;
			RESULT_337 <= RESULT_P26;
			RESULT_529 <= RESULT_P37;
			RESULT_689 <= RESULT_P48;
			RESULT_80 <= RESULT_P14;
			RESULT_304 <= RESULT_P25;
			RESULT_496 <= RESULT_P36;
			RESULT_656 <= RESULT_P47;
			RESULT_784 <= RESULT_P58;
			RESULT_47 <= RESULT_P13;
			RESULT_271 <= RESULT_P24;
			RESULT_463 <= RESULT_P35;
			RESULT_623 <= RESULT_P46;
			RESULT_751 <= RESULT_P57;
			RESULT_847 <= RESULT_P68;
			RESULT_14 <= RESULT_P12;
			RESULT_238 <= RESULT_P23;
			RESULT_430 <= RESULT_P34;
			RESULT_590 <= RESULT_P45;
			RESULT_718 <= RESULT_P56;
			RESULT_814 <= RESULT_P67;
			RESULT_878 <= RESULT_P78;
			end
			24: begin
			RESULT_213 <= RESULT_P18;
			RESULT_180 <= RESULT_P17;
			RESULT_404 <= RESULT_P28;
			RESULT_147 <= RESULT_P16;
			RESULT_371 <= RESULT_P27;
			RESULT_563 <= RESULT_P38;
			RESULT_114 <= RESULT_P15;
			RESULT_338 <= RESULT_P26;
			RESULT_530 <= RESULT_P37;
			RESULT_690 <= RESULT_P48;
			RESULT_81 <= RESULT_P14;
			RESULT_305 <= RESULT_P25;
			RESULT_497 <= RESULT_P36;
			RESULT_657 <= RESULT_P47;
			RESULT_785 <= RESULT_P58;
			RESULT_48 <= RESULT_P13;
			RESULT_272 <= RESULT_P24;
			RESULT_464 <= RESULT_P35;
			RESULT_624 <= RESULT_P46;
			RESULT_752 <= RESULT_P57;
			RESULT_848 <= RESULT_P68;
			RESULT_15 <= RESULT_P12;
			RESULT_239 <= RESULT_P23;
			RESULT_431 <= RESULT_P34;
			RESULT_591 <= RESULT_P45;
			RESULT_719 <= RESULT_P56;
			RESULT_815 <= RESULT_P67;
			RESULT_879 <= RESULT_P78;
			end
			25: begin
			RESULT_214 <= RESULT_P18;
			RESULT_181 <= RESULT_P17;
			RESULT_405 <= RESULT_P28;
			RESULT_148 <= RESULT_P16;
			RESULT_372 <= RESULT_P27;
			RESULT_564 <= RESULT_P38;
			RESULT_115 <= RESULT_P15;
			RESULT_339 <= RESULT_P26;
			RESULT_531 <= RESULT_P37;
			RESULT_691 <= RESULT_P48;
			RESULT_82 <= RESULT_P14;
			RESULT_306 <= RESULT_P25;
			RESULT_498 <= RESULT_P36;
			RESULT_658 <= RESULT_P47;
			RESULT_786 <= RESULT_P58;
			RESULT_49 <= RESULT_P13;
			RESULT_273 <= RESULT_P24;
			RESULT_465 <= RESULT_P35;
			RESULT_625 <= RESULT_P46;
			RESULT_753 <= RESULT_P57;
			RESULT_849 <= RESULT_P68;
			RESULT_16 <= RESULT_P12;
			RESULT_240 <= RESULT_P23;
			RESULT_432 <= RESULT_P34;
			RESULT_592 <= RESULT_P45;
			RESULT_720 <= RESULT_P56;
			RESULT_816 <= RESULT_P67;
			RESULT_880 <= RESULT_P78;
			end
			26: begin
			RESULT_215 <= RESULT_P18;
			RESULT_182 <= RESULT_P17;
			RESULT_406 <= RESULT_P28;
			RESULT_149 <= RESULT_P16;
			RESULT_373 <= RESULT_P27;
			RESULT_565 <= RESULT_P38;
			RESULT_116 <= RESULT_P15;
			RESULT_340 <= RESULT_P26;
			RESULT_532 <= RESULT_P37;
			RESULT_692 <= RESULT_P48;
			RESULT_83 <= RESULT_P14;
			RESULT_307 <= RESULT_P25;
			RESULT_499 <= RESULT_P36;
			RESULT_659 <= RESULT_P47;
			RESULT_787 <= RESULT_P58;
			RESULT_50 <= RESULT_P13;
			RESULT_274 <= RESULT_P24;
			RESULT_466 <= RESULT_P35;
			RESULT_626 <= RESULT_P46;
			RESULT_754 <= RESULT_P57;
			RESULT_850 <= RESULT_P68;
			RESULT_17 <= RESULT_P12;
			RESULT_241 <= RESULT_P23;
			RESULT_433 <= RESULT_P34;
			RESULT_593 <= RESULT_P45;
			RESULT_721 <= RESULT_P56;
			RESULT_817 <= RESULT_P67;
			RESULT_881 <= RESULT_P78;
			end
			27: begin
			RESULT_216 <= RESULT_P18;
			RESULT_183 <= RESULT_P17;
			RESULT_407 <= RESULT_P28;
			RESULT_150 <= RESULT_P16;
			RESULT_374 <= RESULT_P27;
			RESULT_566 <= RESULT_P38;
			RESULT_117 <= RESULT_P15;
			RESULT_341 <= RESULT_P26;
			RESULT_533 <= RESULT_P37;
			RESULT_693 <= RESULT_P48;
			RESULT_84 <= RESULT_P14;
			RESULT_308 <= RESULT_P25;
			RESULT_500 <= RESULT_P36;
			RESULT_660 <= RESULT_P47;
			RESULT_788 <= RESULT_P58;
			RESULT_51 <= RESULT_P13;
			RESULT_275 <= RESULT_P24;
			RESULT_467 <= RESULT_P35;
			RESULT_627 <= RESULT_P46;
			RESULT_755 <= RESULT_P57;
			RESULT_851 <= RESULT_P68;
			RESULT_18 <= RESULT_P12;
			RESULT_242 <= RESULT_P23;
			RESULT_434 <= RESULT_P34;
			RESULT_594 <= RESULT_P45;
			RESULT_722 <= RESULT_P56;
			RESULT_818 <= RESULT_P67;
			RESULT_882 <= RESULT_P78;
			end
			28: begin
			RESULT_217 <= RESULT_P18;
			RESULT_184 <= RESULT_P17;
			RESULT_408 <= RESULT_P28;
			RESULT_151 <= RESULT_P16;
			RESULT_375 <= RESULT_P27;
			RESULT_567 <= RESULT_P38;
			RESULT_118 <= RESULT_P15;
			RESULT_342 <= RESULT_P26;
			RESULT_534 <= RESULT_P37;
			RESULT_694 <= RESULT_P48;
			RESULT_85 <= RESULT_P14;
			RESULT_309 <= RESULT_P25;
			RESULT_501 <= RESULT_P36;
			RESULT_661 <= RESULT_P47;
			RESULT_789 <= RESULT_P58;
			RESULT_52 <= RESULT_P13;
			RESULT_276 <= RESULT_P24;
			RESULT_468 <= RESULT_P35;
			RESULT_628 <= RESULT_P46;
			RESULT_756 <= RESULT_P57;
			RESULT_852 <= RESULT_P68;
			RESULT_19 <= RESULT_P12;
			RESULT_243 <= RESULT_P23;
			RESULT_435 <= RESULT_P34;
			RESULT_595 <= RESULT_P45;
			RESULT_723 <= RESULT_P56;
			RESULT_819 <= RESULT_P67;
			RESULT_883 <= RESULT_P78;
			end
			29: begin
			RESULT_218 <= RESULT_P18;
			RESULT_185 <= RESULT_P17;
			RESULT_409 <= RESULT_P28;
			RESULT_152 <= RESULT_P16;
			RESULT_376 <= RESULT_P27;
			RESULT_568 <= RESULT_P38;
			RESULT_119 <= RESULT_P15;
			RESULT_343 <= RESULT_P26;
			RESULT_535 <= RESULT_P37;
			RESULT_695 <= RESULT_P48;
			RESULT_86 <= RESULT_P14;
			RESULT_310 <= RESULT_P25;
			RESULT_502 <= RESULT_P36;
			RESULT_662 <= RESULT_P47;
			RESULT_790 <= RESULT_P58;
			RESULT_53 <= RESULT_P13;
			RESULT_277 <= RESULT_P24;
			RESULT_469 <= RESULT_P35;
			RESULT_629 <= RESULT_P46;
			RESULT_757 <= RESULT_P57;
			RESULT_853 <= RESULT_P68;
			RESULT_20 <= RESULT_P12;
			RESULT_244 <= RESULT_P23;
			RESULT_436 <= RESULT_P34;
			RESULT_596 <= RESULT_P45;
			RESULT_724 <= RESULT_P56;
			RESULT_820 <= RESULT_P67;
			RESULT_884 <= RESULT_P78;
			end
			30: begin
			RESULT_219 <= RESULT_P18;
			RESULT_186 <= RESULT_P17;
			RESULT_410 <= RESULT_P28;
			RESULT_153 <= RESULT_P16;
			RESULT_377 <= RESULT_P27;
			RESULT_569 <= RESULT_P38;
			RESULT_120 <= RESULT_P15;
			RESULT_344 <= RESULT_P26;
			RESULT_536 <= RESULT_P37;
			RESULT_696 <= RESULT_P48;
			RESULT_87 <= RESULT_P14;
			RESULT_311 <= RESULT_P25;
			RESULT_503 <= RESULT_P36;
			RESULT_663 <= RESULT_P47;
			RESULT_791 <= RESULT_P58;
			RESULT_54 <= RESULT_P13;
			RESULT_278 <= RESULT_P24;
			RESULT_470 <= RESULT_P35;
			RESULT_630 <= RESULT_P46;
			RESULT_758 <= RESULT_P57;
			RESULT_854 <= RESULT_P68;
			RESULT_21 <= RESULT_P12;
			RESULT_245 <= RESULT_P23;
			RESULT_437 <= RESULT_P34;
			RESULT_597 <= RESULT_P45;
			RESULT_725 <= RESULT_P56;
			RESULT_821 <= RESULT_P67;
			RESULT_885 <= RESULT_P78;
			end
			31: begin
			RESULT_220 <= RESULT_P18;
			RESULT_187 <= RESULT_P17;
			RESULT_411 <= RESULT_P28;
			RESULT_154 <= RESULT_P16;
			RESULT_378 <= RESULT_P27;
			RESULT_570 <= RESULT_P38;
			RESULT_121 <= RESULT_P15;
			RESULT_345 <= RESULT_P26;
			RESULT_537 <= RESULT_P37;
			RESULT_697 <= RESULT_P48;
			RESULT_88 <= RESULT_P14;
			RESULT_312 <= RESULT_P25;
			RESULT_504 <= RESULT_P36;
			RESULT_664 <= RESULT_P47;
			RESULT_792 <= RESULT_P58;
			RESULT_55 <= RESULT_P13;
			RESULT_279 <= RESULT_P24;
			RESULT_471 <= RESULT_P35;
			RESULT_631 <= RESULT_P46;
			RESULT_759 <= RESULT_P57;
			RESULT_855 <= RESULT_P68;
			RESULT_22 <= RESULT_P12;
			RESULT_246 <= RESULT_P23;
			RESULT_438 <= RESULT_P34;
			RESULT_598 <= RESULT_P45;
			RESULT_726 <= RESULT_P56;
			RESULT_822 <= RESULT_P67;
			RESULT_886 <= RESULT_P78;
			end
			32: begin
			RESULT_221 <= RESULT_P18;
			RESULT_188 <= RESULT_P17;
			RESULT_412 <= RESULT_P28;
			RESULT_155 <= RESULT_P16;
			RESULT_379 <= RESULT_P27;
			RESULT_571 <= RESULT_P38;
			RESULT_122 <= RESULT_P15;
			RESULT_346 <= RESULT_P26;
			RESULT_538 <= RESULT_P37;
			RESULT_698 <= RESULT_P48;
			RESULT_89 <= RESULT_P14;
			RESULT_313 <= RESULT_P25;
			RESULT_505 <= RESULT_P36;
			RESULT_665 <= RESULT_P47;
			RESULT_793 <= RESULT_P58;
			RESULT_56 <= RESULT_P13;
			RESULT_280 <= RESULT_P24;
			RESULT_472 <= RESULT_P35;
			RESULT_632 <= RESULT_P46;
			RESULT_760 <= RESULT_P57;
			RESULT_856 <= RESULT_P68;
			RESULT_23 <= RESULT_P12;
			RESULT_247 <= RESULT_P23;
			RESULT_439 <= RESULT_P34;
			RESULT_599 <= RESULT_P45;
			RESULT_727 <= RESULT_P56;
			RESULT_823 <= RESULT_P67;
			RESULT_887 <= RESULT_P78;
			end
			33: begin
			RESULT_222 <= RESULT_P18;
			RESULT_189 <= RESULT_P17;
			RESULT_413 <= RESULT_P28;
			RESULT_156 <= RESULT_P16;
			RESULT_380 <= RESULT_P27;
			RESULT_572 <= RESULT_P38;
			RESULT_123 <= RESULT_P15;
			RESULT_347 <= RESULT_P26;
			RESULT_539 <= RESULT_P37;
			RESULT_699 <= RESULT_P48;
			RESULT_90 <= RESULT_P14;
			RESULT_314 <= RESULT_P25;
			RESULT_506 <= RESULT_P36;
			RESULT_666 <= RESULT_P47;
			RESULT_794 <= RESULT_P58;
			RESULT_57 <= RESULT_P13;
			RESULT_281 <= RESULT_P24;
			RESULT_473 <= RESULT_P35;
			RESULT_633 <= RESULT_P46;
			RESULT_761 <= RESULT_P57;
			RESULT_857 <= RESULT_P68;
			RESULT_24 <= RESULT_P12;
			RESULT_248 <= RESULT_P23;
			RESULT_440 <= RESULT_P34;
			RESULT_600 <= RESULT_P45;
			RESULT_728 <= RESULT_P56;
			RESULT_824 <= RESULT_P67;
			RESULT_888 <= RESULT_P78;
			end
			34: begin
			RESULT_223 <= RESULT_P18;
			RESULT_190 <= RESULT_P17;
			RESULT_414 <= RESULT_P28;
			RESULT_157 <= RESULT_P16;
			RESULT_381 <= RESULT_P27;
			RESULT_573 <= RESULT_P38;
			RESULT_124 <= RESULT_P15;
			RESULT_348 <= RESULT_P26;
			RESULT_540 <= RESULT_P37;
			RESULT_700 <= RESULT_P48;
			RESULT_91 <= RESULT_P14;
			RESULT_315 <= RESULT_P25;
			RESULT_507 <= RESULT_P36;
			RESULT_667 <= RESULT_P47;
			RESULT_795 <= RESULT_P58;
			RESULT_58 <= RESULT_P13;
			RESULT_282 <= RESULT_P24;
			RESULT_474 <= RESULT_P35;
			RESULT_634 <= RESULT_P46;
			RESULT_762 <= RESULT_P57;
			RESULT_858 <= RESULT_P68;
			RESULT_25 <= RESULT_P12;
			RESULT_249 <= RESULT_P23;
			RESULT_441 <= RESULT_P34;
			RESULT_601 <= RESULT_P45;
			RESULT_729 <= RESULT_P56;
			RESULT_825 <= RESULT_P67;
			RESULT_889 <= RESULT_P78;
			end
			35: begin
			RESULT_191 <= RESULT_P17;
			RESULT_415 <= RESULT_P28;
			RESULT_158 <= RESULT_P16;
			RESULT_382 <= RESULT_P27;
			RESULT_574 <= RESULT_P38;
			RESULT_125 <= RESULT_P15;
			RESULT_349 <= RESULT_P26;
			RESULT_541 <= RESULT_P37;
			RESULT_701 <= RESULT_P48;
			RESULT_92 <= RESULT_P14;
			RESULT_316 <= RESULT_P25;
			RESULT_508 <= RESULT_P36;
			RESULT_668 <= RESULT_P47;
			RESULT_796 <= RESULT_P58;
			RESULT_59 <= RESULT_P13;
			RESULT_283 <= RESULT_P24;
			RESULT_475 <= RESULT_P35;
			RESULT_635 <= RESULT_P46;
			RESULT_763 <= RESULT_P57;
			RESULT_859 <= RESULT_P68;
			RESULT_26 <= RESULT_P12;
			RESULT_250 <= RESULT_P23;
			RESULT_442 <= RESULT_P34;
			RESULT_602 <= RESULT_P45;
			RESULT_730 <= RESULT_P56;
			RESULT_826 <= RESULT_P67;
			RESULT_890 <= RESULT_P78;
			end
			36: begin
			RESULT_159 <= RESULT_P16;
			RESULT_383 <= RESULT_P27;
			RESULT_575 <= RESULT_P38;
			RESULT_126 <= RESULT_P15;
			RESULT_350 <= RESULT_P26;
			RESULT_542 <= RESULT_P37;
			RESULT_702 <= RESULT_P48;
			RESULT_93 <= RESULT_P14;
			RESULT_317 <= RESULT_P25;
			RESULT_509 <= RESULT_P36;
			RESULT_669 <= RESULT_P47;
			RESULT_797 <= RESULT_P58;
			RESULT_60 <= RESULT_P13;
			RESULT_284 <= RESULT_P24;
			RESULT_476 <= RESULT_P35;
			RESULT_636 <= RESULT_P46;
			RESULT_764 <= RESULT_P57;
			RESULT_860 <= RESULT_P68;
			RESULT_27 <= RESULT_P12;
			RESULT_251 <= RESULT_P23;
			RESULT_443 <= RESULT_P34;
			RESULT_603 <= RESULT_P45;
			RESULT_731 <= RESULT_P56;
			RESULT_827 <= RESULT_P67;
			RESULT_891 <= RESULT_P78;
			end
			37: begin
			RESULT_127 <= RESULT_P15;
			RESULT_351 <= RESULT_P26;
			RESULT_543 <= RESULT_P37;
			RESULT_703 <= RESULT_P48;
			RESULT_94 <= RESULT_P14;
			RESULT_318 <= RESULT_P25;
			RESULT_510 <= RESULT_P36;
			RESULT_670 <= RESULT_P47;
			RESULT_798 <= RESULT_P58;
			RESULT_61 <= RESULT_P13;
			RESULT_285 <= RESULT_P24;
			RESULT_477 <= RESULT_P35;
			RESULT_637 <= RESULT_P46;
			RESULT_765 <= RESULT_P57;
			RESULT_861 <= RESULT_P68;
			RESULT_28 <= RESULT_P12;
			RESULT_252 <= RESULT_P23;
			RESULT_444 <= RESULT_P34;
			RESULT_604 <= RESULT_P45;
			RESULT_732 <= RESULT_P56;
			RESULT_828 <= RESULT_P67;
			RESULT_892 <= RESULT_P78;
			end
			38: begin
			RESULT_95 <= RESULT_P14;
			RESULT_319 <= RESULT_P25;
			RESULT_511 <= RESULT_P36;
			RESULT_671 <= RESULT_P47;
			RESULT_799 <= RESULT_P58;
			RESULT_62 <= RESULT_P13;
			RESULT_286 <= RESULT_P24;
			RESULT_478 <= RESULT_P35;
			RESULT_638 <= RESULT_P46;
			RESULT_766 <= RESULT_P57;
			RESULT_862 <= RESULT_P68;
			RESULT_29 <= RESULT_P12;
			RESULT_253 <= RESULT_P23;
			RESULT_445 <= RESULT_P34;
			RESULT_605 <= RESULT_P45;
			RESULT_733 <= RESULT_P56;
			RESULT_829 <= RESULT_P67;
			RESULT_893 <= RESULT_P78;
			end
			39: begin
			RESULT_63 <= RESULT_P13;
			RESULT_287 <= RESULT_P24;
			RESULT_479 <= RESULT_P35;
			RESULT_639 <= RESULT_P46;
			RESULT_767 <= RESULT_P57;
			RESULT_863 <= RESULT_P68;
			RESULT_30 <= RESULT_P12;
			RESULT_254 <= RESULT_P23;
			RESULT_446 <= RESULT_P34;
			RESULT_606 <= RESULT_P45;
			RESULT_734 <= RESULT_P56;
			RESULT_830 <= RESULT_P67;
			RESULT_894 <= RESULT_P78;
			end
			40: begin
			RESULT_31 <= RESULT_P12;
			RESULT_255 <= RESULT_P23;
			RESULT_447 <= RESULT_P34;
			RESULT_607 <= RESULT_P45;
			RESULT_735 <= RESULT_P56;
			RESULT_831 <= RESULT_P67;
			RESULT_895 <= RESULT_P78;
			end

            default: begin
                 RESULT_0 <= 16'b0;
				 RESULT_1 <= 16'b0;
				 RESULT_2 <= 16'b0;
				 RESULT_3 <= 16'b0;
				 RESULT_4 <= 16'b0;
				 RESULT_5 <= 16'b0;
				 RESULT_6 <= 16'b0;
				 RESULT_7 <= 16'b0;
				 RESULT_8 <= 16'b0;
				 RESULT_9 <= 16'b0;
				 RESULT_10 <= 16'b0;
				 RESULT_11 <= 16'b0;
				 RESULT_12 <= 16'b0;
				 RESULT_13 <= 16'b0;
				 RESULT_14 <= 16'b0;
				 RESULT_15 <= 16'b0;
				 RESULT_16 <= 16'b0;
				 RESULT_17 <= 16'b0;
				 RESULT_18 <= 16'b0;
				 RESULT_19 <= 16'b0;
				 RESULT_20 <= 16'b0;
				 RESULT_21 <= 16'b0;
				 RESULT_22 <= 16'b0;
				 RESULT_23 <= 16'b0;
				 RESULT_24 <= 16'b0;
				 RESULT_25 <= 16'b0;
				 RESULT_26 <= 16'b0;
				 RESULT_27 <= 16'b0;
				 RESULT_28 <= 16'b0;
				 RESULT_29 <= 16'b0;
				 RESULT_30 <= 16'b0;
				 RESULT_31 <= 16'b0;
				 RESULT_32 <= 16'b0;
				 RESULT_33 <= 16'b0;
				 RESULT_34 <= 16'b0;
				 RESULT_35 <= 16'b0;
				 RESULT_36 <= 16'b0;
				 RESULT_37 <= 16'b0;
				 RESULT_38 <= 16'b0;
				 RESULT_39 <= 16'b0;
				 RESULT_40 <= 16'b0;
				 RESULT_41 <= 16'b0;
				 RESULT_42 <= 16'b0;
				 RESULT_43 <= 16'b0;
				 RESULT_44 <= 16'b0;
				 RESULT_45 <= 16'b0;
				 RESULT_46 <= 16'b0;
				 RESULT_47 <= 16'b0;
				 RESULT_48 <= 16'b0;
				 RESULT_49 <= 16'b0;
				 RESULT_50 <= 16'b0;
				 RESULT_51 <= 16'b0;
				 RESULT_52 <= 16'b0;
				 RESULT_53 <= 16'b0;
				 RESULT_54 <= 16'b0;
				 RESULT_55 <= 16'b0;
				 RESULT_56 <= 16'b0;
				 RESULT_57 <= 16'b0;
				 RESULT_58 <= 16'b0;
				 RESULT_59 <= 16'b0;
				 RESULT_60 <= 16'b0;
				 RESULT_61 <= 16'b0;
				 RESULT_62 <= 16'b0;
				 RESULT_63 <= 16'b0;
				 RESULT_64 <= 16'b0;
				 RESULT_65 <= 16'b0;
				 RESULT_66 <= 16'b0;
				 RESULT_67 <= 16'b0;
				 RESULT_68 <= 16'b0;
				 RESULT_69 <= 16'b0;
				 RESULT_70 <= 16'b0;
				 RESULT_71 <= 16'b0;
				 RESULT_72 <= 16'b0;
				 RESULT_73 <= 16'b0;
				 RESULT_74 <= 16'b0;
				 RESULT_75 <= 16'b0;
				 RESULT_76 <= 16'b0;
				 RESULT_77 <= 16'b0;
				 RESULT_78 <= 16'b0;
				 RESULT_79 <= 16'b0;
				 RESULT_80 <= 16'b0;
				 RESULT_81 <= 16'b0;
				 RESULT_82 <= 16'b0;
				 RESULT_83 <= 16'b0;
				 RESULT_84 <= 16'b0;
				 RESULT_85 <= 16'b0;
				 RESULT_86 <= 16'b0;
				 RESULT_87 <= 16'b0;
				 RESULT_88 <= 16'b0;
				 RESULT_89 <= 16'b0;
				 RESULT_90 <= 16'b0;
				 RESULT_91 <= 16'b0;
				 RESULT_92 <= 16'b0;
				 RESULT_93 <= 16'b0;
				 RESULT_94 <= 16'b0;
				 RESULT_95 <= 16'b0;
				 RESULT_96 <= 16'b0;
				 RESULT_97 <= 16'b0;
				 RESULT_98 <= 16'b0;
				 RESULT_99 <= 16'b0;
				 RESULT_100 <= 16'b0;
				 RESULT_101 <= 16'b0;
				 RESULT_102 <= 16'b0;
				 RESULT_103 <= 16'b0;
				 RESULT_104 <= 16'b0;
				 RESULT_105 <= 16'b0;
				 RESULT_106 <= 16'b0;
				 RESULT_107 <= 16'b0;
				 RESULT_108 <= 16'b0;
				 RESULT_109 <= 16'b0;
				 RESULT_110 <= 16'b0;
				 RESULT_111 <= 16'b0;
				 RESULT_112 <= 16'b0;
				 RESULT_113 <= 16'b0;
				 RESULT_114 <= 16'b0;
				 RESULT_115 <= 16'b0;
				 RESULT_116 <= 16'b0;
				 RESULT_117 <= 16'b0;
				 RESULT_118 <= 16'b0;
				 RESULT_119 <= 16'b0;
				 RESULT_120 <= 16'b0;
				 RESULT_121 <= 16'b0;
				 RESULT_122 <= 16'b0;
				 RESULT_123 <= 16'b0;
				 RESULT_124 <= 16'b0;
				 RESULT_125 <= 16'b0;
				 RESULT_126 <= 16'b0;
				 RESULT_127 <= 16'b0;
				 RESULT_128 <= 16'b0;
				 RESULT_129 <= 16'b0;
				 RESULT_130 <= 16'b0;
				 RESULT_131 <= 16'b0;
				 RESULT_132 <= 16'b0;
				 RESULT_133 <= 16'b0;
				 RESULT_134 <= 16'b0;
				 RESULT_135 <= 16'b0;
				 RESULT_136 <= 16'b0;
				 RESULT_137 <= 16'b0;
				 RESULT_138 <= 16'b0;
				 RESULT_139 <= 16'b0;
				 RESULT_140 <= 16'b0;
				 RESULT_141 <= 16'b0;
				 RESULT_142 <= 16'b0;
				 RESULT_143 <= 16'b0;
				 RESULT_144 <= 16'b0;
				 RESULT_145 <= 16'b0;
				 RESULT_146 <= 16'b0;
				 RESULT_147 <= 16'b0;
				 RESULT_148 <= 16'b0;
				 RESULT_149 <= 16'b0;
				 RESULT_150 <= 16'b0;
				 RESULT_151 <= 16'b0;
				 RESULT_152 <= 16'b0;
				 RESULT_153 <= 16'b0;
				 RESULT_154 <= 16'b0;
				 RESULT_155 <= 16'b0;
				 RESULT_156 <= 16'b0;
				 RESULT_157 <= 16'b0;
				 RESULT_158 <= 16'b0;
				 RESULT_159 <= 16'b0;
				 RESULT_160 <= 16'b0;
				 RESULT_161 <= 16'b0;
				 RESULT_162 <= 16'b0;
				 RESULT_163 <= 16'b0;
				 RESULT_164 <= 16'b0;
				 RESULT_165 <= 16'b0;
				 RESULT_166 <= 16'b0;
				 RESULT_167 <= 16'b0;
				 RESULT_168 <= 16'b0;
				 RESULT_169 <= 16'b0;
				 RESULT_170 <= 16'b0;
				 RESULT_171 <= 16'b0;
				 RESULT_172 <= 16'b0;
				 RESULT_173 <= 16'b0;
				 RESULT_174 <= 16'b0;
				 RESULT_175 <= 16'b0;
				 RESULT_176 <= 16'b0;
				 RESULT_177 <= 16'b0;
				 RESULT_178 <= 16'b0;
				 RESULT_179 <= 16'b0;
				 RESULT_180 <= 16'b0;
				 RESULT_181 <= 16'b0;
				 RESULT_182 <= 16'b0;
				 RESULT_183 <= 16'b0;
				 RESULT_184 <= 16'b0;
				 RESULT_185 <= 16'b0;
				 RESULT_186 <= 16'b0;
				 RESULT_187 <= 16'b0;
				 RESULT_188 <= 16'b0;
				 RESULT_189 <= 16'b0;
				 RESULT_190 <= 16'b0;
				 RESULT_191 <= 16'b0;
				 RESULT_192 <= 16'b0;
				 RESULT_193 <= 16'b0;
				 RESULT_194 <= 16'b0;
				 RESULT_195 <= 16'b0;
				 RESULT_196 <= 16'b0;
				 RESULT_197 <= 16'b0;
				 RESULT_198 <= 16'b0;
				 RESULT_199 <= 16'b0;
				 RESULT_200 <= 16'b0;
				 RESULT_201 <= 16'b0;
				 RESULT_202 <= 16'b0;
				 RESULT_203 <= 16'b0;
				 RESULT_204 <= 16'b0;
				 RESULT_205 <= 16'b0;
				 RESULT_206 <= 16'b0;
				 RESULT_207 <= 16'b0;
				 RESULT_208 <= 16'b0;
				 RESULT_209 <= 16'b0;
				 RESULT_210 <= 16'b0;
				 RESULT_211 <= 16'b0;
				 RESULT_212 <= 16'b0;
				 RESULT_213 <= 16'b0;
				 RESULT_214 <= 16'b0;
				 RESULT_215 <= 16'b0;
				 RESULT_216 <= 16'b0;
				 RESULT_217 <= 16'b0;
				 RESULT_218 <= 16'b0;
				 RESULT_219 <= 16'b0;
				 RESULT_220 <= 16'b0;
				 RESULT_221 <= 16'b0;
				 RESULT_222 <= 16'b0;
				 RESULT_223 <= 16'b0;
				 RESULT_224 <= 16'b0;
				 RESULT_225 <= 16'b0;
				 RESULT_226 <= 16'b0;
				 RESULT_227 <= 16'b0;
				 RESULT_228 <= 16'b0;
				 RESULT_229 <= 16'b0;
				 RESULT_230 <= 16'b0;
				 RESULT_231 <= 16'b0;
				 RESULT_232 <= 16'b0;
				 RESULT_233 <= 16'b0;
				 RESULT_234 <= 16'b0;
				 RESULT_235 <= 16'b0;
				 RESULT_236 <= 16'b0;
				 RESULT_237 <= 16'b0;
				 RESULT_238 <= 16'b0;
				 RESULT_239 <= 16'b0;
				 RESULT_240 <= 16'b0;
				 RESULT_241 <= 16'b0;
				 RESULT_242 <= 16'b0;
				 RESULT_243 <= 16'b0;
				 RESULT_244 <= 16'b0;
				 RESULT_245 <= 16'b0;
				 RESULT_246 <= 16'b0;
				 RESULT_247 <= 16'b0;
				 RESULT_248 <= 16'b0;
				 RESULT_249 <= 16'b0;
				 RESULT_250 <= 16'b0;
				 RESULT_251 <= 16'b0;
				 RESULT_252 <= 16'b0;
				 RESULT_253 <= 16'b0;
				 RESULT_254 <= 16'b0;
				 RESULT_255 <= 16'b0;
				 RESULT_256 <= 16'b0;
				 RESULT_257 <= 16'b0;
				 RESULT_258 <= 16'b0;
				 RESULT_259 <= 16'b0;
				 RESULT_260 <= 16'b0;
				 RESULT_261 <= 16'b0;
				 RESULT_262 <= 16'b0;
				 RESULT_263 <= 16'b0;
				 RESULT_264 <= 16'b0;
				 RESULT_265 <= 16'b0;
				 RESULT_266 <= 16'b0;
				 RESULT_267 <= 16'b0;
				 RESULT_268 <= 16'b0;
				 RESULT_269 <= 16'b0;
				 RESULT_270 <= 16'b0;
				 RESULT_271 <= 16'b0;
				 RESULT_272 <= 16'b0;
				 RESULT_273 <= 16'b0;
				 RESULT_274 <= 16'b0;
				 RESULT_275 <= 16'b0;
				 RESULT_276 <= 16'b0;
				 RESULT_277 <= 16'b0;
				 RESULT_278 <= 16'b0;
				 RESULT_279 <= 16'b0;
				 RESULT_280 <= 16'b0;
				 RESULT_281 <= 16'b0;
				 RESULT_282 <= 16'b0;
				 RESULT_283 <= 16'b0;
				 RESULT_284 <= 16'b0;
				 RESULT_285 <= 16'b0;
				 RESULT_286 <= 16'b0;
				 RESULT_287 <= 16'b0;
				 RESULT_288 <= 16'b0;
				 RESULT_289 <= 16'b0;
				 RESULT_290 <= 16'b0;
				 RESULT_291 <= 16'b0;
				 RESULT_292 <= 16'b0;
				 RESULT_293 <= 16'b0;
				 RESULT_294 <= 16'b0;
				 RESULT_295 <= 16'b0;
				 RESULT_296 <= 16'b0;
				 RESULT_297 <= 16'b0;
				 RESULT_298 <= 16'b0;
				 RESULT_299 <= 16'b0;
				 RESULT_300 <= 16'b0;
				 RESULT_301 <= 16'b0;
				 RESULT_302 <= 16'b0;
				 RESULT_303 <= 16'b0;
				 RESULT_304 <= 16'b0;
				 RESULT_305 <= 16'b0;
				 RESULT_306 <= 16'b0;
				 RESULT_307 <= 16'b0;
				 RESULT_308 <= 16'b0;
				 RESULT_309 <= 16'b0;
				 RESULT_310 <= 16'b0;
				 RESULT_311 <= 16'b0;
				 RESULT_312 <= 16'b0;
				 RESULT_313 <= 16'b0;
				 RESULT_314 <= 16'b0;
				 RESULT_315 <= 16'b0;
				 RESULT_316 <= 16'b0;
				 RESULT_317 <= 16'b0;
				 RESULT_318 <= 16'b0;
				 RESULT_319 <= 16'b0;
				 RESULT_320 <= 16'b0;
				 RESULT_321 <= 16'b0;
				 RESULT_322 <= 16'b0;
				 RESULT_323 <= 16'b0;
				 RESULT_324 <= 16'b0;
				 RESULT_325 <= 16'b0;
				 RESULT_326 <= 16'b0;
				 RESULT_327 <= 16'b0;
				 RESULT_328 <= 16'b0;
				 RESULT_329 <= 16'b0;
				 RESULT_330 <= 16'b0;
				 RESULT_331 <= 16'b0;
				 RESULT_332 <= 16'b0;
				 RESULT_333 <= 16'b0;
				 RESULT_334 <= 16'b0;
				 RESULT_335 <= 16'b0;
				 RESULT_336 <= 16'b0;
				 RESULT_337 <= 16'b0;
				 RESULT_338 <= 16'b0;
				 RESULT_339 <= 16'b0;
				 RESULT_340 <= 16'b0;
				 RESULT_341 <= 16'b0;
				 RESULT_342 <= 16'b0;
				 RESULT_343 <= 16'b0;
				 RESULT_344 <= 16'b0;
				 RESULT_345 <= 16'b0;
				 RESULT_346 <= 16'b0;
				 RESULT_347 <= 16'b0;
				 RESULT_348 <= 16'b0;
				 RESULT_349 <= 16'b0;
				 RESULT_350 <= 16'b0;
				 RESULT_351 <= 16'b0;
				 RESULT_352 <= 16'b0;
				 RESULT_353 <= 16'b0;
				 RESULT_354 <= 16'b0;
				 RESULT_355 <= 16'b0;
				 RESULT_356 <= 16'b0;
				 RESULT_357 <= 16'b0;
				 RESULT_358 <= 16'b0;
				 RESULT_359 <= 16'b0;
				 RESULT_360 <= 16'b0;
				 RESULT_361 <= 16'b0;
				 RESULT_362 <= 16'b0;
				 RESULT_363 <= 16'b0;
				 RESULT_364 <= 16'b0;
				 RESULT_365 <= 16'b0;
				 RESULT_366 <= 16'b0;
				 RESULT_367 <= 16'b0;
				 RESULT_368 <= 16'b0;
				 RESULT_369 <= 16'b0;
				 RESULT_370 <= 16'b0;
				 RESULT_371 <= 16'b0;
				 RESULT_372 <= 16'b0;
				 RESULT_373 <= 16'b0;
				 RESULT_374 <= 16'b0;
				 RESULT_375 <= 16'b0;
				 RESULT_376 <= 16'b0;
				 RESULT_377 <= 16'b0;
				 RESULT_378 <= 16'b0;
				 RESULT_379 <= 16'b0;
				 RESULT_380 <= 16'b0;
				 RESULT_381 <= 16'b0;
				 RESULT_382 <= 16'b0;
				 RESULT_383 <= 16'b0;
				 RESULT_384 <= 16'b0;
				 RESULT_385 <= 16'b0;
				 RESULT_386 <= 16'b0;
				 RESULT_387 <= 16'b0;
				 RESULT_388 <= 16'b0;
				 RESULT_389 <= 16'b0;
				 RESULT_390 <= 16'b0;
				 RESULT_391 <= 16'b0;
				 RESULT_392 <= 16'b0;
				 RESULT_393 <= 16'b0;
				 RESULT_394 <= 16'b0;
				 RESULT_395 <= 16'b0;
				 RESULT_396 <= 16'b0;
				 RESULT_397 <= 16'b0;
				 RESULT_398 <= 16'b0;
				 RESULT_399 <= 16'b0;
				 RESULT_400 <= 16'b0;
				 RESULT_401 <= 16'b0;
				 RESULT_402 <= 16'b0;
				 RESULT_403 <= 16'b0;
				 RESULT_404 <= 16'b0;
				 RESULT_405 <= 16'b0;
				 RESULT_406 <= 16'b0;
				 RESULT_407 <= 16'b0;
				 RESULT_408 <= 16'b0;
				 RESULT_409 <= 16'b0;
				 RESULT_410 <= 16'b0;
				 RESULT_411 <= 16'b0;
				 RESULT_412 <= 16'b0;
				 RESULT_413 <= 16'b0;
				 RESULT_414 <= 16'b0;
				 RESULT_415 <= 16'b0;
				 RESULT_416 <= 16'b0;
				 RESULT_417 <= 16'b0;
				 RESULT_418 <= 16'b0;
				 RESULT_419 <= 16'b0;
				 RESULT_420 <= 16'b0;
				 RESULT_421 <= 16'b0;
				 RESULT_422 <= 16'b0;
				 RESULT_423 <= 16'b0;
				 RESULT_424 <= 16'b0;
				 RESULT_425 <= 16'b0;
				 RESULT_426 <= 16'b0;
				 RESULT_427 <= 16'b0;
				 RESULT_428 <= 16'b0;
				 RESULT_429 <= 16'b0;
				 RESULT_430 <= 16'b0;
				 RESULT_431 <= 16'b0;
				 RESULT_432 <= 16'b0;
				 RESULT_433 <= 16'b0;
				 RESULT_434 <= 16'b0;
				 RESULT_435 <= 16'b0;
				 RESULT_436 <= 16'b0;
				 RESULT_437 <= 16'b0;
				 RESULT_438 <= 16'b0;
				 RESULT_439 <= 16'b0;
				 RESULT_440 <= 16'b0;
				 RESULT_441 <= 16'b0;
				 RESULT_442 <= 16'b0;
				 RESULT_443 <= 16'b0;
				 RESULT_444 <= 16'b0;
				 RESULT_445 <= 16'b0;
				 RESULT_446 <= 16'b0;
				 RESULT_447 <= 16'b0;
				 RESULT_448 <= 16'b0;
				 RESULT_449 <= 16'b0;
				 RESULT_450 <= 16'b0;
				 RESULT_451 <= 16'b0;
				 RESULT_452 <= 16'b0;
				 RESULT_453 <= 16'b0;
				 RESULT_454 <= 16'b0;
				 RESULT_455 <= 16'b0;
				 RESULT_456 <= 16'b0;
				 RESULT_457 <= 16'b0;
				 RESULT_458 <= 16'b0;
				 RESULT_459 <= 16'b0;
				 RESULT_460 <= 16'b0;
				 RESULT_461 <= 16'b0;
				 RESULT_462 <= 16'b0;
				 RESULT_463 <= 16'b0;
				 RESULT_464 <= 16'b0;
				 RESULT_465 <= 16'b0;
				 RESULT_466 <= 16'b0;
				 RESULT_467 <= 16'b0;
				 RESULT_468 <= 16'b0;
				 RESULT_469 <= 16'b0;
				 RESULT_470 <= 16'b0;
				 RESULT_471 <= 16'b0;
				 RESULT_472 <= 16'b0;
				 RESULT_473 <= 16'b0;
				 RESULT_474 <= 16'b0;
				 RESULT_475 <= 16'b0;
				 RESULT_476 <= 16'b0;
				 RESULT_477 <= 16'b0;
				 RESULT_478 <= 16'b0;
				 RESULT_479 <= 16'b0;
				 RESULT_480 <= 16'b0;
				 RESULT_481 <= 16'b0;
				 RESULT_482 <= 16'b0;
				 RESULT_483 <= 16'b0;
				 RESULT_484 <= 16'b0;
				 RESULT_485 <= 16'b0;
				 RESULT_486 <= 16'b0;
				 RESULT_487 <= 16'b0;
				 RESULT_488 <= 16'b0;
				 RESULT_489 <= 16'b0;
				 RESULT_490 <= 16'b0;
				 RESULT_491 <= 16'b0;
				 RESULT_492 <= 16'b0;
				 RESULT_493 <= 16'b0;
				 RESULT_494 <= 16'b0;
				 RESULT_495 <= 16'b0;
				 RESULT_496 <= 16'b0;
				 RESULT_497 <= 16'b0;
				 RESULT_498 <= 16'b0;
				 RESULT_499 <= 16'b0;
				 RESULT_500 <= 16'b0;
				 RESULT_501 <= 16'b0;
				 RESULT_502 <= 16'b0;
				 RESULT_503 <= 16'b0;
				 RESULT_504 <= 16'b0;
				 RESULT_505 <= 16'b0;
				 RESULT_506 <= 16'b0;
				 RESULT_507 <= 16'b0;
				 RESULT_508 <= 16'b0;
				 RESULT_509 <= 16'b0;
				 RESULT_510 <= 16'b0;
				 RESULT_511 <= 16'b0;
				 RESULT_512 <= 16'b0;
				 RESULT_513 <= 16'b0;
				 RESULT_514 <= 16'b0;
				 RESULT_515 <= 16'b0;
				 RESULT_516 <= 16'b0;
				 RESULT_517 <= 16'b0;
				 RESULT_518 <= 16'b0;
				 RESULT_519 <= 16'b0;
				 RESULT_520 <= 16'b0;
				 RESULT_521 <= 16'b0;
				 RESULT_522 <= 16'b0;
				 RESULT_523 <= 16'b0;
				 RESULT_524 <= 16'b0;
				 RESULT_525 <= 16'b0;
				 RESULT_526 <= 16'b0;
				 RESULT_527 <= 16'b0;
				 RESULT_528 <= 16'b0;
				 RESULT_529 <= 16'b0;
				 RESULT_530 <= 16'b0;
				 RESULT_531 <= 16'b0;
				 RESULT_532 <= 16'b0;
				 RESULT_533 <= 16'b0;
				 RESULT_534 <= 16'b0;
				 RESULT_535 <= 16'b0;
				 RESULT_536 <= 16'b0;
				 RESULT_537 <= 16'b0;
				 RESULT_538 <= 16'b0;
				 RESULT_539 <= 16'b0;
				 RESULT_540 <= 16'b0;
				 RESULT_541 <= 16'b0;
				 RESULT_542 <= 16'b0;
				 RESULT_543 <= 16'b0;
				 RESULT_544 <= 16'b0;
				 RESULT_545 <= 16'b0;
				 RESULT_546 <= 16'b0;
				 RESULT_547 <= 16'b0;
				 RESULT_548 <= 16'b0;
				 RESULT_549 <= 16'b0;
				 RESULT_550 <= 16'b0;
				 RESULT_551 <= 16'b0;
				 RESULT_552 <= 16'b0;
				 RESULT_553 <= 16'b0;
				 RESULT_554 <= 16'b0;
				 RESULT_555 <= 16'b0;
				 RESULT_556 <= 16'b0;
				 RESULT_557 <= 16'b0;
				 RESULT_558 <= 16'b0;
				 RESULT_559 <= 16'b0;
				 RESULT_560 <= 16'b0;
				 RESULT_561 <= 16'b0;
				 RESULT_562 <= 16'b0;
				 RESULT_563 <= 16'b0;
				 RESULT_564 <= 16'b0;
				 RESULT_565 <= 16'b0;
				 RESULT_566 <= 16'b0;
				 RESULT_567 <= 16'b0;
				 RESULT_568 <= 16'b0;
				 RESULT_569 <= 16'b0;
				 RESULT_570 <= 16'b0;
				 RESULT_571 <= 16'b0;
				 RESULT_572 <= 16'b0;
				 RESULT_573 <= 16'b0;
				 RESULT_574 <= 16'b0;
				 RESULT_575 <= 16'b0;
				 RESULT_576 <= 16'b0;
				 RESULT_577 <= 16'b0;
				 RESULT_578 <= 16'b0;
				 RESULT_579 <= 16'b0;
				 RESULT_580 <= 16'b0;
				 RESULT_581 <= 16'b0;
				 RESULT_582 <= 16'b0;
				 RESULT_583 <= 16'b0;
				 RESULT_584 <= 16'b0;
				 RESULT_585 <= 16'b0;
				 RESULT_586 <= 16'b0;
				 RESULT_587 <= 16'b0;
				 RESULT_588 <= 16'b0;
				 RESULT_589 <= 16'b0;
				 RESULT_590 <= 16'b0;
				 RESULT_591 <= 16'b0;
				 RESULT_592 <= 16'b0;
				 RESULT_593 <= 16'b0;
				 RESULT_594 <= 16'b0;
				 RESULT_595 <= 16'b0;
				 RESULT_596 <= 16'b0;
				 RESULT_597 <= 16'b0;
				 RESULT_598 <= 16'b0;
				 RESULT_599 <= 16'b0;
				 RESULT_600 <= 16'b0;
				 RESULT_601 <= 16'b0;
				 RESULT_602 <= 16'b0;
				 RESULT_603 <= 16'b0;
				 RESULT_604 <= 16'b0;
				 RESULT_605 <= 16'b0;
				 RESULT_606 <= 16'b0;
				 RESULT_607 <= 16'b0;
				 RESULT_608 <= 16'b0;
				 RESULT_609 <= 16'b0;
				 RESULT_610 <= 16'b0;
				 RESULT_611 <= 16'b0;
				 RESULT_612 <= 16'b0;
				 RESULT_613 <= 16'b0;
				 RESULT_614 <= 16'b0;
				 RESULT_615 <= 16'b0;
				 RESULT_616 <= 16'b0;
				 RESULT_617 <= 16'b0;
				 RESULT_618 <= 16'b0;
				 RESULT_619 <= 16'b0;
				 RESULT_620 <= 16'b0;
				 RESULT_621 <= 16'b0;
				 RESULT_622 <= 16'b0;
				 RESULT_623 <= 16'b0;
				 RESULT_624 <= 16'b0;
				 RESULT_625 <= 16'b0;
				 RESULT_626 <= 16'b0;
				 RESULT_627 <= 16'b0;
				 RESULT_628 <= 16'b0;
				 RESULT_629 <= 16'b0;
				 RESULT_630 <= 16'b0;
				 RESULT_631 <= 16'b0;
				 RESULT_632 <= 16'b0;
				 RESULT_633 <= 16'b0;
				 RESULT_634 <= 16'b0;
				 RESULT_635 <= 16'b0;
				 RESULT_636 <= 16'b0;
				 RESULT_637 <= 16'b0;
				 RESULT_638 <= 16'b0;
				 RESULT_639 <= 16'b0;
				 RESULT_640 <= 16'b0;
				 RESULT_641 <= 16'b0;
				 RESULT_642 <= 16'b0;
				 RESULT_643 <= 16'b0;
				 RESULT_644 <= 16'b0;
				 RESULT_645 <= 16'b0;
				 RESULT_646 <= 16'b0;
				 RESULT_647 <= 16'b0;
				 RESULT_648 <= 16'b0;
				 RESULT_649 <= 16'b0;
				 RESULT_650 <= 16'b0;
				 RESULT_651 <= 16'b0;
				 RESULT_652 <= 16'b0;
				 RESULT_653 <= 16'b0;
				 RESULT_654 <= 16'b0;
				 RESULT_655 <= 16'b0;
				 RESULT_656 <= 16'b0;
				 RESULT_657 <= 16'b0;
				 RESULT_658 <= 16'b0;
				 RESULT_659 <= 16'b0;
				 RESULT_660 <= 16'b0;
				 RESULT_661 <= 16'b0;
				 RESULT_662 <= 16'b0;
				 RESULT_663 <= 16'b0;
				 RESULT_664 <= 16'b0;
				 RESULT_665 <= 16'b0;
				 RESULT_666 <= 16'b0;
				 RESULT_667 <= 16'b0;
				 RESULT_668 <= 16'b0;
				 RESULT_669 <= 16'b0;
				 RESULT_670 <= 16'b0;
				 RESULT_671 <= 16'b0;
				 RESULT_672 <= 16'b0;
				 RESULT_673 <= 16'b0;
				 RESULT_674 <= 16'b0;
				 RESULT_675 <= 16'b0;
				 RESULT_676 <= 16'b0;
				 RESULT_677 <= 16'b0;
				 RESULT_678 <= 16'b0;
				 RESULT_679 <= 16'b0;
				 RESULT_680 <= 16'b0;
				 RESULT_681 <= 16'b0;
				 RESULT_682 <= 16'b0;
				 RESULT_683 <= 16'b0;
				 RESULT_684 <= 16'b0;
				 RESULT_685 <= 16'b0;
				 RESULT_686 <= 16'b0;
				 RESULT_687 <= 16'b0;
				 RESULT_688 <= 16'b0;
				 RESULT_689 <= 16'b0;
				 RESULT_690 <= 16'b0;
				 RESULT_691 <= 16'b0;
				 RESULT_692 <= 16'b0;
				 RESULT_693 <= 16'b0;
				 RESULT_694 <= 16'b0;
				 RESULT_695 <= 16'b0;
				 RESULT_696 <= 16'b0;
				 RESULT_697 <= 16'b0;
				 RESULT_698 <= 16'b0;
				 RESULT_699 <= 16'b0;
				 RESULT_700 <= 16'b0;
				 RESULT_701 <= 16'b0;
				 RESULT_702 <= 16'b0;
				 RESULT_703 <= 16'b0;
				 RESULT_704 <= 16'b0;
				 RESULT_705 <= 16'b0;
				 RESULT_706 <= 16'b0;
				 RESULT_707 <= 16'b0;
				 RESULT_708 <= 16'b0;
				 RESULT_709 <= 16'b0;
				 RESULT_710 <= 16'b0;
				 RESULT_711 <= 16'b0;
				 RESULT_712 <= 16'b0;
				 RESULT_713 <= 16'b0;
				 RESULT_714 <= 16'b0;
				 RESULT_715 <= 16'b0;
				 RESULT_716 <= 16'b0;
				 RESULT_717 <= 16'b0;
				 RESULT_718 <= 16'b0;
				 RESULT_719 <= 16'b0;
				 RESULT_720 <= 16'b0;
				 RESULT_721 <= 16'b0;
				 RESULT_722 <= 16'b0;
				 RESULT_723 <= 16'b0;
				 RESULT_724 <= 16'b0;
				 RESULT_725 <= 16'b0;
				 RESULT_726 <= 16'b0;
				 RESULT_727 <= 16'b0;
				 RESULT_728 <= 16'b0;
				 RESULT_729 <= 16'b0;
				 RESULT_730 <= 16'b0;
				 RESULT_731 <= 16'b0;
				 RESULT_732 <= 16'b0;
				 RESULT_733 <= 16'b0;
				 RESULT_734 <= 16'b0;
				 RESULT_735 <= 16'b0;
				 RESULT_736 <= 16'b0;
				 RESULT_737 <= 16'b0;
				 RESULT_738 <= 16'b0;
				 RESULT_739 <= 16'b0;
				 RESULT_740 <= 16'b0;
				 RESULT_741 <= 16'b0;
				 RESULT_742 <= 16'b0;
				 RESULT_743 <= 16'b0;
				 RESULT_744 <= 16'b0;
				 RESULT_745 <= 16'b0;
				 RESULT_746 <= 16'b0;
				 RESULT_747 <= 16'b0;
				 RESULT_748 <= 16'b0;
				 RESULT_749 <= 16'b0;
				 RESULT_750 <= 16'b0;
				 RESULT_751 <= 16'b0;
				 RESULT_752 <= 16'b0;
				 RESULT_753 <= 16'b0;
				 RESULT_754 <= 16'b0;
				 RESULT_755 <= 16'b0;
				 RESULT_756 <= 16'b0;
				 RESULT_757 <= 16'b0;
				 RESULT_758 <= 16'b0;
				 RESULT_759 <= 16'b0;
				 RESULT_760 <= 16'b0;
				 RESULT_761 <= 16'b0;
				 RESULT_762 <= 16'b0;
				 RESULT_763 <= 16'b0;
				 RESULT_764 <= 16'b0;
				 RESULT_765 <= 16'b0;
				 RESULT_766 <= 16'b0;
				 RESULT_767 <= 16'b0;
				 RESULT_768 <= 16'b0;
				 RESULT_769 <= 16'b0;
				 RESULT_770 <= 16'b0;
				 RESULT_771 <= 16'b0;
				 RESULT_772 <= 16'b0;
				 RESULT_773 <= 16'b0;
				 RESULT_774 <= 16'b0;
				 RESULT_775 <= 16'b0;
				 RESULT_776 <= 16'b0;
				 RESULT_777 <= 16'b0;
				 RESULT_778 <= 16'b0;
				 RESULT_779 <= 16'b0;
				 RESULT_780 <= 16'b0;
				 RESULT_781 <= 16'b0;
				 RESULT_782 <= 16'b0;
				 RESULT_783 <= 16'b0;
				 RESULT_784 <= 16'b0;
				 RESULT_785 <= 16'b0;
				 RESULT_786 <= 16'b0;
				 RESULT_787 <= 16'b0;
				 RESULT_788 <= 16'b0;
				 RESULT_789 <= 16'b0;
				 RESULT_790 <= 16'b0;
				 RESULT_791 <= 16'b0;
				 RESULT_792 <= 16'b0;
				 RESULT_793 <= 16'b0;
				 RESULT_794 <= 16'b0;
				 RESULT_795 <= 16'b0;
				 RESULT_796 <= 16'b0;
				 RESULT_797 <= 16'b0;
				 RESULT_798 <= 16'b0;
				 RESULT_799 <= 16'b0;
				 RESULT_800 <= 16'b0;
				 RESULT_801 <= 16'b0;
				 RESULT_802 <= 16'b0;
				 RESULT_803 <= 16'b0;
				 RESULT_804 <= 16'b0;
				 RESULT_805 <= 16'b0;
				 RESULT_806 <= 16'b0;
				 RESULT_807 <= 16'b0;
				 RESULT_808 <= 16'b0;
				 RESULT_809 <= 16'b0;
				 RESULT_810 <= 16'b0;
				 RESULT_811 <= 16'b0;
				 RESULT_812 <= 16'b0;
				 RESULT_813 <= 16'b0;
				 RESULT_814 <= 16'b0;
				 RESULT_815 <= 16'b0;
				 RESULT_816 <= 16'b0;
				 RESULT_817 <= 16'b0;
				 RESULT_818 <= 16'b0;
				 RESULT_819 <= 16'b0;
				 RESULT_820 <= 16'b0;
				 RESULT_821 <= 16'b0;
				 RESULT_822 <= 16'b0;
				 RESULT_823 <= 16'b0;
				 RESULT_824 <= 16'b0;
				 RESULT_825 <= 16'b0;
				 RESULT_826 <= 16'b0;
				 RESULT_827 <= 16'b0;
				 RESULT_828 <= 16'b0;
				 RESULT_829 <= 16'b0;
				 RESULT_830 <= 16'b0;
				 RESULT_831 <= 16'b0;
				 RESULT_832 <= 16'b0;
				 RESULT_833 <= 16'b0;
				 RESULT_834 <= 16'b0;
				 RESULT_835 <= 16'b0;
				 RESULT_836 <= 16'b0;
				 RESULT_837 <= 16'b0;
				 RESULT_838 <= 16'b0;
				 RESULT_839 <= 16'b0;
				 RESULT_840 <= 16'b0;
				 RESULT_841 <= 16'b0;
				 RESULT_842 <= 16'b0;
				 RESULT_843 <= 16'b0;
				 RESULT_844 <= 16'b0;
				 RESULT_845 <= 16'b0;
				 RESULT_846 <= 16'b0;
				 RESULT_847 <= 16'b0;
				 RESULT_848 <= 16'b0;
				 RESULT_849 <= 16'b0;
				 RESULT_850 <= 16'b0;
				 RESULT_851 <= 16'b0;
				 RESULT_852 <= 16'b0;
				 RESULT_853 <= 16'b0;
				 RESULT_854 <= 16'b0;
				 RESULT_855 <= 16'b0;
				 RESULT_856 <= 16'b0;
				 RESULT_857 <= 16'b0;
				 RESULT_858 <= 16'b0;
				 RESULT_859 <= 16'b0;
				 RESULT_860 <= 16'b0;
				 RESULT_861 <= 16'b0;
				 RESULT_862 <= 16'b0;
				 RESULT_863 <= 16'b0;
				 RESULT_864 <= 16'b0;
				 RESULT_865 <= 16'b0;
				 RESULT_866 <= 16'b0;
				 RESULT_867 <= 16'b0;
				 RESULT_868 <= 16'b0;
				 RESULT_869 <= 16'b0;
				 RESULT_870 <= 16'b0;
				 RESULT_871 <= 16'b0;
				 RESULT_872 <= 16'b0;
				 RESULT_873 <= 16'b0;
				 RESULT_874 <= 16'b0;
				 RESULT_875 <= 16'b0;
				 RESULT_876 <= 16'b0;
				 RESULT_877 <= 16'b0;
				 RESULT_878 <= 16'b0;
				 RESULT_879 <= 16'b0;
				 RESULT_880 <= 16'b0;
				 RESULT_881 <= 16'b0;
				 RESULT_882 <= 16'b0;
				 RESULT_883 <= 16'b0;
				 RESULT_884 <= 16'b0;
				 RESULT_885 <= 16'b0;
				 RESULT_886 <= 16'b0;
				 RESULT_887 <= 16'b0;
				 RESULT_888 <= 16'b0;
				 RESULT_889 <= 16'b0;
				 RESULT_890 <= 16'b0;
				 RESULT_891 <= 16'b0;
				 RESULT_892 <= 16'b0;
				 RESULT_893 <= 16'b0;
				 RESULT_894 <= 16'b0;
				 RESULT_895 <= 16'b0;
            end
         endcase
	  end else begin
		RESULT_0 <= 16'b0;
         RESULT_1 <= 16'b0;
         RESULT_2 <= 16'b0;
         RESULT_3 <= 16'b0;
         RESULT_4 <= 16'b0;
         RESULT_5 <= 16'b0;
         RESULT_6 <= 16'b0;
         RESULT_7 <= 16'b0;
         RESULT_8 <= 16'b0;
         RESULT_9 <= 16'b0;
         RESULT_10 <= 16'b0;
         RESULT_11 <= 16'b0;
         RESULT_12 <= 16'b0;
         RESULT_13 <= 16'b0;
         RESULT_14 <= 16'b0;
         RESULT_15 <= 16'b0;
         RESULT_16 <= 16'b0;
         RESULT_17 <= 16'b0;
         RESULT_18 <= 16'b0;
         RESULT_19 <= 16'b0;
         RESULT_20 <= 16'b0;
         RESULT_21 <= 16'b0;
         RESULT_22 <= 16'b0;
         RESULT_23 <= 16'b0;
         RESULT_24 <= 16'b0;
         RESULT_25 <= 16'b0;
         RESULT_26 <= 16'b0;
         RESULT_27 <= 16'b0;
         RESULT_28 <= 16'b0;
         RESULT_29 <= 16'b0;
         RESULT_30 <= 16'b0;
         RESULT_31 <= 16'b0;
         RESULT_32 <= 16'b0;
         RESULT_33 <= 16'b0;
         RESULT_34 <= 16'b0;
         RESULT_35 <= 16'b0;
         RESULT_36 <= 16'b0;
         RESULT_37 <= 16'b0;
         RESULT_38 <= 16'b0;
         RESULT_39 <= 16'b0;
         RESULT_40 <= 16'b0;
         RESULT_41 <= 16'b0;
         RESULT_42 <= 16'b0;
         RESULT_43 <= 16'b0;
         RESULT_44 <= 16'b0;
         RESULT_45 <= 16'b0;
         RESULT_46 <= 16'b0;
         RESULT_47 <= 16'b0;
         RESULT_48 <= 16'b0;
         RESULT_49 <= 16'b0;
         RESULT_50 <= 16'b0;
         RESULT_51 <= 16'b0;
         RESULT_52 <= 16'b0;
         RESULT_53 <= 16'b0;
         RESULT_54 <= 16'b0;
         RESULT_55 <= 16'b0;
         RESULT_56 <= 16'b0;
         RESULT_57 <= 16'b0;
         RESULT_58 <= 16'b0;
         RESULT_59 <= 16'b0;
         RESULT_60 <= 16'b0;
         RESULT_61 <= 16'b0;
         RESULT_62 <= 16'b0;
         RESULT_63 <= 16'b0;
         RESULT_64 <= 16'b0;
         RESULT_65 <= 16'b0;
         RESULT_66 <= 16'b0;
         RESULT_67 <= 16'b0;
         RESULT_68 <= 16'b0;
         RESULT_69 <= 16'b0;
         RESULT_70 <= 16'b0;
         RESULT_71 <= 16'b0;
         RESULT_72 <= 16'b0;
         RESULT_73 <= 16'b0;
         RESULT_74 <= 16'b0;
         RESULT_75 <= 16'b0;
         RESULT_76 <= 16'b0;
         RESULT_77 <= 16'b0;
         RESULT_78 <= 16'b0;
         RESULT_79 <= 16'b0;
         RESULT_80 <= 16'b0;
         RESULT_81 <= 16'b0;
         RESULT_82 <= 16'b0;
         RESULT_83 <= 16'b0;
         RESULT_84 <= 16'b0;
         RESULT_85 <= 16'b0;
         RESULT_86 <= 16'b0;
         RESULT_87 <= 16'b0;
         RESULT_88 <= 16'b0;
         RESULT_89 <= 16'b0;
         RESULT_90 <= 16'b0;
         RESULT_91 <= 16'b0;
         RESULT_92 <= 16'b0;
         RESULT_93 <= 16'b0;
         RESULT_94 <= 16'b0;
         RESULT_95 <= 16'b0;
         RESULT_96 <= 16'b0;
         RESULT_97 <= 16'b0;
         RESULT_98 <= 16'b0;
         RESULT_99 <= 16'b0;
         RESULT_100 <= 16'b0;
         RESULT_101 <= 16'b0;
         RESULT_102 <= 16'b0;
         RESULT_103 <= 16'b0;
         RESULT_104 <= 16'b0;
         RESULT_105 <= 16'b0;
         RESULT_106 <= 16'b0;
         RESULT_107 <= 16'b0;
         RESULT_108 <= 16'b0;
         RESULT_109 <= 16'b0;
         RESULT_110 <= 16'b0;
         RESULT_111 <= 16'b0;
         RESULT_112 <= 16'b0;
         RESULT_113 <= 16'b0;
         RESULT_114 <= 16'b0;
         RESULT_115 <= 16'b0;
         RESULT_116 <= 16'b0;
         RESULT_117 <= 16'b0;
         RESULT_118 <= 16'b0;
         RESULT_119 <= 16'b0;
         RESULT_120 <= 16'b0;
         RESULT_121 <= 16'b0;
         RESULT_122 <= 16'b0;
         RESULT_123 <= 16'b0;
         RESULT_124 <= 16'b0;
         RESULT_125 <= 16'b0;
         RESULT_126 <= 16'b0;
         RESULT_127 <= 16'b0;
         RESULT_128 <= 16'b0;
         RESULT_129 <= 16'b0;
         RESULT_130 <= 16'b0;
         RESULT_131 <= 16'b0;
         RESULT_132 <= 16'b0;
         RESULT_133 <= 16'b0;
         RESULT_134 <= 16'b0;
         RESULT_135 <= 16'b0;
         RESULT_136 <= 16'b0;
         RESULT_137 <= 16'b0;
         RESULT_138 <= 16'b0;
         RESULT_139 <= 16'b0;
         RESULT_140 <= 16'b0;
         RESULT_141 <= 16'b0;
         RESULT_142 <= 16'b0;
         RESULT_143 <= 16'b0;
         RESULT_144 <= 16'b0;
         RESULT_145 <= 16'b0;
         RESULT_146 <= 16'b0;
         RESULT_147 <= 16'b0;
         RESULT_148 <= 16'b0;
         RESULT_149 <= 16'b0;
         RESULT_150 <= 16'b0;
         RESULT_151 <= 16'b0;
         RESULT_152 <= 16'b0;
         RESULT_153 <= 16'b0;
         RESULT_154 <= 16'b0;
         RESULT_155 <= 16'b0;
         RESULT_156 <= 16'b0;
         RESULT_157 <= 16'b0;
         RESULT_158 <= 16'b0;
         RESULT_159 <= 16'b0;
         RESULT_160 <= 16'b0;
         RESULT_161 <= 16'b0;
         RESULT_162 <= 16'b0;
         RESULT_163 <= 16'b0;
         RESULT_164 <= 16'b0;
         RESULT_165 <= 16'b0;
         RESULT_166 <= 16'b0;
         RESULT_167 <= 16'b0;
         RESULT_168 <= 16'b0;
         RESULT_169 <= 16'b0;
         RESULT_170 <= 16'b0;
         RESULT_171 <= 16'b0;
         RESULT_172 <= 16'b0;
         RESULT_173 <= 16'b0;
         RESULT_174 <= 16'b0;
         RESULT_175 <= 16'b0;
         RESULT_176 <= 16'b0;
         RESULT_177 <= 16'b0;
         RESULT_178 <= 16'b0;
         RESULT_179 <= 16'b0;
         RESULT_180 <= 16'b0;
         RESULT_181 <= 16'b0;
         RESULT_182 <= 16'b0;
         RESULT_183 <= 16'b0;
         RESULT_184 <= 16'b0;
         RESULT_185 <= 16'b0;
         RESULT_186 <= 16'b0;
         RESULT_187 <= 16'b0;
         RESULT_188 <= 16'b0;
         RESULT_189 <= 16'b0;
         RESULT_190 <= 16'b0;
         RESULT_191 <= 16'b0;
         RESULT_192 <= 16'b0;
         RESULT_193 <= 16'b0;
         RESULT_194 <= 16'b0;
         RESULT_195 <= 16'b0;
         RESULT_196 <= 16'b0;
         RESULT_197 <= 16'b0;
         RESULT_198 <= 16'b0;
         RESULT_199 <= 16'b0;
         RESULT_200 <= 16'b0;
         RESULT_201 <= 16'b0;
         RESULT_202 <= 16'b0;
         RESULT_203 <= 16'b0;
         RESULT_204 <= 16'b0;
         RESULT_205 <= 16'b0;
         RESULT_206 <= 16'b0;
         RESULT_207 <= 16'b0;
         RESULT_208 <= 16'b0;
         RESULT_209 <= 16'b0;
         RESULT_210 <= 16'b0;
         RESULT_211 <= 16'b0;
         RESULT_212 <= 16'b0;
         RESULT_213 <= 16'b0;
         RESULT_214 <= 16'b0;
         RESULT_215 <= 16'b0;
         RESULT_216 <= 16'b0;
         RESULT_217 <= 16'b0;
         RESULT_218 <= 16'b0;
         RESULT_219 <= 16'b0;
         RESULT_220 <= 16'b0;
         RESULT_221 <= 16'b0;
         RESULT_222 <= 16'b0;
         RESULT_223 <= 16'b0;
         RESULT_224 <= 16'b0;
         RESULT_225 <= 16'b0;
         RESULT_226 <= 16'b0;
         RESULT_227 <= 16'b0;
         RESULT_228 <= 16'b0;
         RESULT_229 <= 16'b0;
         RESULT_230 <= 16'b0;
         RESULT_231 <= 16'b0;
         RESULT_232 <= 16'b0;
         RESULT_233 <= 16'b0;
         RESULT_234 <= 16'b0;
         RESULT_235 <= 16'b0;
         RESULT_236 <= 16'b0;
         RESULT_237 <= 16'b0;
         RESULT_238 <= 16'b0;
         RESULT_239 <= 16'b0;
         RESULT_240 <= 16'b0;
         RESULT_241 <= 16'b0;
         RESULT_242 <= 16'b0;
         RESULT_243 <= 16'b0;
         RESULT_244 <= 16'b0;
         RESULT_245 <= 16'b0;
         RESULT_246 <= 16'b0;
         RESULT_247 <= 16'b0;
         RESULT_248 <= 16'b0;
         RESULT_249 <= 16'b0;
         RESULT_250 <= 16'b0;
         RESULT_251 <= 16'b0;
         RESULT_252 <= 16'b0;
         RESULT_253 <= 16'b0;
         RESULT_254 <= 16'b0;
         RESULT_255 <= 16'b0;
         RESULT_256 <= 16'b0;
         RESULT_257 <= 16'b0;
         RESULT_258 <= 16'b0;
         RESULT_259 <= 16'b0;
         RESULT_260 <= 16'b0;
         RESULT_261 <= 16'b0;
         RESULT_262 <= 16'b0;
         RESULT_263 <= 16'b0;
         RESULT_264 <= 16'b0;
         RESULT_265 <= 16'b0;
         RESULT_266 <= 16'b0;
         RESULT_267 <= 16'b0;
         RESULT_268 <= 16'b0;
         RESULT_269 <= 16'b0;
         RESULT_270 <= 16'b0;
         RESULT_271 <= 16'b0;
         RESULT_272 <= 16'b0;
         RESULT_273 <= 16'b0;
         RESULT_274 <= 16'b0;
         RESULT_275 <= 16'b0;
         RESULT_276 <= 16'b0;
         RESULT_277 <= 16'b0;
         RESULT_278 <= 16'b0;
         RESULT_279 <= 16'b0;
         RESULT_280 <= 16'b0;
         RESULT_281 <= 16'b0;
         RESULT_282 <= 16'b0;
         RESULT_283 <= 16'b0;
         RESULT_284 <= 16'b0;
         RESULT_285 <= 16'b0;
         RESULT_286 <= 16'b0;
         RESULT_287 <= 16'b0;
         RESULT_288 <= 16'b0;
         RESULT_289 <= 16'b0;
         RESULT_290 <= 16'b0;
         RESULT_291 <= 16'b0;
         RESULT_292 <= 16'b0;
         RESULT_293 <= 16'b0;
         RESULT_294 <= 16'b0;
         RESULT_295 <= 16'b0;
         RESULT_296 <= 16'b0;
         RESULT_297 <= 16'b0;
         RESULT_298 <= 16'b0;
         RESULT_299 <= 16'b0;
         RESULT_300 <= 16'b0;
         RESULT_301 <= 16'b0;
         RESULT_302 <= 16'b0;
         RESULT_303 <= 16'b0;
         RESULT_304 <= 16'b0;
         RESULT_305 <= 16'b0;
         RESULT_306 <= 16'b0;
         RESULT_307 <= 16'b0;
         RESULT_308 <= 16'b0;
         RESULT_309 <= 16'b0;
         RESULT_310 <= 16'b0;
         RESULT_311 <= 16'b0;
         RESULT_312 <= 16'b0;
         RESULT_313 <= 16'b0;
         RESULT_314 <= 16'b0;
         RESULT_315 <= 16'b0;
         RESULT_316 <= 16'b0;
         RESULT_317 <= 16'b0;
         RESULT_318 <= 16'b0;
         RESULT_319 <= 16'b0;
         RESULT_320 <= 16'b0;
         RESULT_321 <= 16'b0;
         RESULT_322 <= 16'b0;
         RESULT_323 <= 16'b0;
         RESULT_324 <= 16'b0;
         RESULT_325 <= 16'b0;
         RESULT_326 <= 16'b0;
         RESULT_327 <= 16'b0;
         RESULT_328 <= 16'b0;
         RESULT_329 <= 16'b0;
         RESULT_330 <= 16'b0;
         RESULT_331 <= 16'b0;
         RESULT_332 <= 16'b0;
         RESULT_333 <= 16'b0;
         RESULT_334 <= 16'b0;
         RESULT_335 <= 16'b0;
         RESULT_336 <= 16'b0;
         RESULT_337 <= 16'b0;
         RESULT_338 <= 16'b0;
         RESULT_339 <= 16'b0;
         RESULT_340 <= 16'b0;
         RESULT_341 <= 16'b0;
         RESULT_342 <= 16'b0;
         RESULT_343 <= 16'b0;
         RESULT_344 <= 16'b0;
         RESULT_345 <= 16'b0;
         RESULT_346 <= 16'b0;
         RESULT_347 <= 16'b0;
         RESULT_348 <= 16'b0;
         RESULT_349 <= 16'b0;
         RESULT_350 <= 16'b0;
         RESULT_351 <= 16'b0;
         RESULT_352 <= 16'b0;
         RESULT_353 <= 16'b0;
         RESULT_354 <= 16'b0;
         RESULT_355 <= 16'b0;
         RESULT_356 <= 16'b0;
         RESULT_357 <= 16'b0;
         RESULT_358 <= 16'b0;
         RESULT_359 <= 16'b0;
         RESULT_360 <= 16'b0;
         RESULT_361 <= 16'b0;
         RESULT_362 <= 16'b0;
         RESULT_363 <= 16'b0;
         RESULT_364 <= 16'b0;
         RESULT_365 <= 16'b0;
         RESULT_366 <= 16'b0;
         RESULT_367 <= 16'b0;
         RESULT_368 <= 16'b0;
         RESULT_369 <= 16'b0;
         RESULT_370 <= 16'b0;
         RESULT_371 <= 16'b0;
         RESULT_372 <= 16'b0;
         RESULT_373 <= 16'b0;
         RESULT_374 <= 16'b0;
         RESULT_375 <= 16'b0;
         RESULT_376 <= 16'b0;
         RESULT_377 <= 16'b0;
         RESULT_378 <= 16'b0;
         RESULT_379 <= 16'b0;
         RESULT_380 <= 16'b0;
         RESULT_381 <= 16'b0;
         RESULT_382 <= 16'b0;
         RESULT_383 <= 16'b0;
         RESULT_384 <= 16'b0;
         RESULT_385 <= 16'b0;
         RESULT_386 <= 16'b0;
         RESULT_387 <= 16'b0;
         RESULT_388 <= 16'b0;
         RESULT_389 <= 16'b0;
         RESULT_390 <= 16'b0;
         RESULT_391 <= 16'b0;
         RESULT_392 <= 16'b0;
         RESULT_393 <= 16'b0;
         RESULT_394 <= 16'b0;
         RESULT_395 <= 16'b0;
         RESULT_396 <= 16'b0;
         RESULT_397 <= 16'b0;
         RESULT_398 <= 16'b0;
         RESULT_399 <= 16'b0;
         RESULT_400 <= 16'b0;
         RESULT_401 <= 16'b0;
         RESULT_402 <= 16'b0;
         RESULT_403 <= 16'b0;
         RESULT_404 <= 16'b0;
         RESULT_405 <= 16'b0;
         RESULT_406 <= 16'b0;
         RESULT_407 <= 16'b0;
         RESULT_408 <= 16'b0;
         RESULT_409 <= 16'b0;
         RESULT_410 <= 16'b0;
         RESULT_411 <= 16'b0;
         RESULT_412 <= 16'b0;
         RESULT_413 <= 16'b0;
         RESULT_414 <= 16'b0;
         RESULT_415 <= 16'b0;
         RESULT_416 <= 16'b0;
         RESULT_417 <= 16'b0;
         RESULT_418 <= 16'b0;
         RESULT_419 <= 16'b0;
         RESULT_420 <= 16'b0;
         RESULT_421 <= 16'b0;
         RESULT_422 <= 16'b0;
         RESULT_423 <= 16'b0;
         RESULT_424 <= 16'b0;
         RESULT_425 <= 16'b0;
         RESULT_426 <= 16'b0;
         RESULT_427 <= 16'b0;
         RESULT_428 <= 16'b0;
         RESULT_429 <= 16'b0;
         RESULT_430 <= 16'b0;
         RESULT_431 <= 16'b0;
         RESULT_432 <= 16'b0;
         RESULT_433 <= 16'b0;
         RESULT_434 <= 16'b0;
         RESULT_435 <= 16'b0;
         RESULT_436 <= 16'b0;
         RESULT_437 <= 16'b0;
         RESULT_438 <= 16'b0;
         RESULT_439 <= 16'b0;
         RESULT_440 <= 16'b0;
         RESULT_441 <= 16'b0;
         RESULT_442 <= 16'b0;
         RESULT_443 <= 16'b0;
         RESULT_444 <= 16'b0;
         RESULT_445 <= 16'b0;
         RESULT_446 <= 16'b0;
         RESULT_447 <= 16'b0;
         RESULT_448 <= 16'b0;
         RESULT_449 <= 16'b0;
         RESULT_450 <= 16'b0;
         RESULT_451 <= 16'b0;
         RESULT_452 <= 16'b0;
         RESULT_453 <= 16'b0;
         RESULT_454 <= 16'b0;
         RESULT_455 <= 16'b0;
         RESULT_456 <= 16'b0;
         RESULT_457 <= 16'b0;
         RESULT_458 <= 16'b0;
         RESULT_459 <= 16'b0;
         RESULT_460 <= 16'b0;
         RESULT_461 <= 16'b0;
         RESULT_462 <= 16'b0;
         RESULT_463 <= 16'b0;
         RESULT_464 <= 16'b0;
         RESULT_465 <= 16'b0;
         RESULT_466 <= 16'b0;
         RESULT_467 <= 16'b0;
         RESULT_468 <= 16'b0;
         RESULT_469 <= 16'b0;
         RESULT_470 <= 16'b0;
         RESULT_471 <= 16'b0;
         RESULT_472 <= 16'b0;
         RESULT_473 <= 16'b0;
         RESULT_474 <= 16'b0;
         RESULT_475 <= 16'b0;
         RESULT_476 <= 16'b0;
         RESULT_477 <= 16'b0;
         RESULT_478 <= 16'b0;
         RESULT_479 <= 16'b0;
         RESULT_480 <= 16'b0;
         RESULT_481 <= 16'b0;
         RESULT_482 <= 16'b0;
         RESULT_483 <= 16'b0;
         RESULT_484 <= 16'b0;
         RESULT_485 <= 16'b0;
         RESULT_486 <= 16'b0;
         RESULT_487 <= 16'b0;
         RESULT_488 <= 16'b0;
         RESULT_489 <= 16'b0;
         RESULT_490 <= 16'b0;
         RESULT_491 <= 16'b0;
         RESULT_492 <= 16'b0;
         RESULT_493 <= 16'b0;
         RESULT_494 <= 16'b0;
         RESULT_495 <= 16'b0;
         RESULT_496 <= 16'b0;
         RESULT_497 <= 16'b0;
         RESULT_498 <= 16'b0;
         RESULT_499 <= 16'b0;
         RESULT_500 <= 16'b0;
         RESULT_501 <= 16'b0;
         RESULT_502 <= 16'b0;
         RESULT_503 <= 16'b0;
         RESULT_504 <= 16'b0;
         RESULT_505 <= 16'b0;
         RESULT_506 <= 16'b0;
         RESULT_507 <= 16'b0;
         RESULT_508 <= 16'b0;
         RESULT_509 <= 16'b0;
         RESULT_510 <= 16'b0;
         RESULT_511 <= 16'b0;
         RESULT_512 <= 16'b0;
         RESULT_513 <= 16'b0;
         RESULT_514 <= 16'b0;
         RESULT_515 <= 16'b0;
         RESULT_516 <= 16'b0;
         RESULT_517 <= 16'b0;
         RESULT_518 <= 16'b0;
         RESULT_519 <= 16'b0;
         RESULT_520 <= 16'b0;
         RESULT_521 <= 16'b0;
         RESULT_522 <= 16'b0;
         RESULT_523 <= 16'b0;
         RESULT_524 <= 16'b0;
         RESULT_525 <= 16'b0;
         RESULT_526 <= 16'b0;
         RESULT_527 <= 16'b0;
         RESULT_528 <= 16'b0;
         RESULT_529 <= 16'b0;
         RESULT_530 <= 16'b0;
         RESULT_531 <= 16'b0;
         RESULT_532 <= 16'b0;
         RESULT_533 <= 16'b0;
         RESULT_534 <= 16'b0;
         RESULT_535 <= 16'b0;
         RESULT_536 <= 16'b0;
         RESULT_537 <= 16'b0;
         RESULT_538 <= 16'b0;
         RESULT_539 <= 16'b0;
         RESULT_540 <= 16'b0;
         RESULT_541 <= 16'b0;
         RESULT_542 <= 16'b0;
         RESULT_543 <= 16'b0;
         RESULT_544 <= 16'b0;
         RESULT_545 <= 16'b0;
         RESULT_546 <= 16'b0;
         RESULT_547 <= 16'b0;
         RESULT_548 <= 16'b0;
         RESULT_549 <= 16'b0;
         RESULT_550 <= 16'b0;
         RESULT_551 <= 16'b0;
         RESULT_552 <= 16'b0;
         RESULT_553 <= 16'b0;
         RESULT_554 <= 16'b0;
         RESULT_555 <= 16'b0;
         RESULT_556 <= 16'b0;
         RESULT_557 <= 16'b0;
         RESULT_558 <= 16'b0;
         RESULT_559 <= 16'b0;
         RESULT_560 <= 16'b0;
         RESULT_561 <= 16'b0;
         RESULT_562 <= 16'b0;
         RESULT_563 <= 16'b0;
         RESULT_564 <= 16'b0;
         RESULT_565 <= 16'b0;
         RESULT_566 <= 16'b0;
         RESULT_567 <= 16'b0;
         RESULT_568 <= 16'b0;
         RESULT_569 <= 16'b0;
         RESULT_570 <= 16'b0;
         RESULT_571 <= 16'b0;
         RESULT_572 <= 16'b0;
         RESULT_573 <= 16'b0;
         RESULT_574 <= 16'b0;
         RESULT_575 <= 16'b0;
         RESULT_576 <= 16'b0;
         RESULT_577 <= 16'b0;
         RESULT_578 <= 16'b0;
         RESULT_579 <= 16'b0;
         RESULT_580 <= 16'b0;
         RESULT_581 <= 16'b0;
         RESULT_582 <= 16'b0;
         RESULT_583 <= 16'b0;
         RESULT_584 <= 16'b0;
         RESULT_585 <= 16'b0;
         RESULT_586 <= 16'b0;
         RESULT_587 <= 16'b0;
         RESULT_588 <= 16'b0;
         RESULT_589 <= 16'b0;
         RESULT_590 <= 16'b0;
         RESULT_591 <= 16'b0;
         RESULT_592 <= 16'b0;
         RESULT_593 <= 16'b0;
         RESULT_594 <= 16'b0;
         RESULT_595 <= 16'b0;
         RESULT_596 <= 16'b0;
         RESULT_597 <= 16'b0;
         RESULT_598 <= 16'b0;
         RESULT_599 <= 16'b0;
         RESULT_600 <= 16'b0;
         RESULT_601 <= 16'b0;
         RESULT_602 <= 16'b0;
         RESULT_603 <= 16'b0;
         RESULT_604 <= 16'b0;
         RESULT_605 <= 16'b0;
         RESULT_606 <= 16'b0;
         RESULT_607 <= 16'b0;
         RESULT_608 <= 16'b0;
         RESULT_609 <= 16'b0;
         RESULT_610 <= 16'b0;
         RESULT_611 <= 16'b0;
         RESULT_612 <= 16'b0;
         RESULT_613 <= 16'b0;
         RESULT_614 <= 16'b0;
         RESULT_615 <= 16'b0;
         RESULT_616 <= 16'b0;
         RESULT_617 <= 16'b0;
         RESULT_618 <= 16'b0;
         RESULT_619 <= 16'b0;
         RESULT_620 <= 16'b0;
         RESULT_621 <= 16'b0;
         RESULT_622 <= 16'b0;
         RESULT_623 <= 16'b0;
         RESULT_624 <= 16'b0;
         RESULT_625 <= 16'b0;
         RESULT_626 <= 16'b0;
         RESULT_627 <= 16'b0;
         RESULT_628 <= 16'b0;
         RESULT_629 <= 16'b0;
         RESULT_630 <= 16'b0;
         RESULT_631 <= 16'b0;
         RESULT_632 <= 16'b0;
         RESULT_633 <= 16'b0;
         RESULT_634 <= 16'b0;
         RESULT_635 <= 16'b0;
         RESULT_636 <= 16'b0;
         RESULT_637 <= 16'b0;
         RESULT_638 <= 16'b0;
         RESULT_639 <= 16'b0;
         RESULT_640 <= 16'b0;
         RESULT_641 <= 16'b0;
         RESULT_642 <= 16'b0;
         RESULT_643 <= 16'b0;
         RESULT_644 <= 16'b0;
         RESULT_645 <= 16'b0;
         RESULT_646 <= 16'b0;
         RESULT_647 <= 16'b0;
         RESULT_648 <= 16'b0;
         RESULT_649 <= 16'b0;
         RESULT_650 <= 16'b0;
         RESULT_651 <= 16'b0;
         RESULT_652 <= 16'b0;
         RESULT_653 <= 16'b0;
         RESULT_654 <= 16'b0;
         RESULT_655 <= 16'b0;
         RESULT_656 <= 16'b0;
         RESULT_657 <= 16'b0;
         RESULT_658 <= 16'b0;
         RESULT_659 <= 16'b0;
         RESULT_660 <= 16'b0;
         RESULT_661 <= 16'b0;
         RESULT_662 <= 16'b0;
         RESULT_663 <= 16'b0;
         RESULT_664 <= 16'b0;
         RESULT_665 <= 16'b0;
         RESULT_666 <= 16'b0;
         RESULT_667 <= 16'b0;
         RESULT_668 <= 16'b0;
         RESULT_669 <= 16'b0;
         RESULT_670 <= 16'b0;
         RESULT_671 <= 16'b0;
         RESULT_672 <= 16'b0;
         RESULT_673 <= 16'b0;
         RESULT_674 <= 16'b0;
         RESULT_675 <= 16'b0;
         RESULT_676 <= 16'b0;
         RESULT_677 <= 16'b0;
         RESULT_678 <= 16'b0;
         RESULT_679 <= 16'b0;
         RESULT_680 <= 16'b0;
         RESULT_681 <= 16'b0;
         RESULT_682 <= 16'b0;
         RESULT_683 <= 16'b0;
         RESULT_684 <= 16'b0;
         RESULT_685 <= 16'b0;
         RESULT_686 <= 16'b0;
         RESULT_687 <= 16'b0;
         RESULT_688 <= 16'b0;
         RESULT_689 <= 16'b0;
         RESULT_690 <= 16'b0;
         RESULT_691 <= 16'b0;
         RESULT_692 <= 16'b0;
         RESULT_693 <= 16'b0;
         RESULT_694 <= 16'b0;
         RESULT_695 <= 16'b0;
         RESULT_696 <= 16'b0;
         RESULT_697 <= 16'b0;
         RESULT_698 <= 16'b0;
         RESULT_699 <= 16'b0;
         RESULT_700 <= 16'b0;
         RESULT_701 <= 16'b0;
         RESULT_702 <= 16'b0;
         RESULT_703 <= 16'b0;
         RESULT_704 <= 16'b0;
         RESULT_705 <= 16'b0;
         RESULT_706 <= 16'b0;
         RESULT_707 <= 16'b0;
         RESULT_708 <= 16'b0;
         RESULT_709 <= 16'b0;
         RESULT_710 <= 16'b0;
         RESULT_711 <= 16'b0;
         RESULT_712 <= 16'b0;
         RESULT_713 <= 16'b0;
         RESULT_714 <= 16'b0;
         RESULT_715 <= 16'b0;
         RESULT_716 <= 16'b0;
         RESULT_717 <= 16'b0;
         RESULT_718 <= 16'b0;
         RESULT_719 <= 16'b0;
         RESULT_720 <= 16'b0;
         RESULT_721 <= 16'b0;
         RESULT_722 <= 16'b0;
         RESULT_723 <= 16'b0;
         RESULT_724 <= 16'b0;
         RESULT_725 <= 16'b0;
         RESULT_726 <= 16'b0;
         RESULT_727 <= 16'b0;
         RESULT_728 <= 16'b0;
         RESULT_729 <= 16'b0;
         RESULT_730 <= 16'b0;
         RESULT_731 <= 16'b0;
         RESULT_732 <= 16'b0;
         RESULT_733 <= 16'b0;
         RESULT_734 <= 16'b0;
         RESULT_735 <= 16'b0;
         RESULT_736 <= 16'b0;
         RESULT_737 <= 16'b0;
         RESULT_738 <= 16'b0;
         RESULT_739 <= 16'b0;
         RESULT_740 <= 16'b0;
         RESULT_741 <= 16'b0;
         RESULT_742 <= 16'b0;
         RESULT_743 <= 16'b0;
         RESULT_744 <= 16'b0;
         RESULT_745 <= 16'b0;
         RESULT_746 <= 16'b0;
         RESULT_747 <= 16'b0;
         RESULT_748 <= 16'b0;
         RESULT_749 <= 16'b0;
         RESULT_750 <= 16'b0;
         RESULT_751 <= 16'b0;
         RESULT_752 <= 16'b0;
         RESULT_753 <= 16'b0;
         RESULT_754 <= 16'b0;
         RESULT_755 <= 16'b0;
         RESULT_756 <= 16'b0;
         RESULT_757 <= 16'b0;
         RESULT_758 <= 16'b0;
         RESULT_759 <= 16'b0;
         RESULT_760 <= 16'b0;
         RESULT_761 <= 16'b0;
         RESULT_762 <= 16'b0;
         RESULT_763 <= 16'b0;
         RESULT_764 <= 16'b0;
         RESULT_765 <= 16'b0;
         RESULT_766 <= 16'b0;
         RESULT_767 <= 16'b0;
         RESULT_768 <= 16'b0;
         RESULT_769 <= 16'b0;
         RESULT_770 <= 16'b0;
         RESULT_771 <= 16'b0;
         RESULT_772 <= 16'b0;
         RESULT_773 <= 16'b0;
         RESULT_774 <= 16'b0;
         RESULT_775 <= 16'b0;
         RESULT_776 <= 16'b0;
         RESULT_777 <= 16'b0;
         RESULT_778 <= 16'b0;
         RESULT_779 <= 16'b0;
         RESULT_780 <= 16'b0;
         RESULT_781 <= 16'b0;
         RESULT_782 <= 16'b0;
         RESULT_783 <= 16'b0;
         RESULT_784 <= 16'b0;
         RESULT_785 <= 16'b0;
         RESULT_786 <= 16'b0;
         RESULT_787 <= 16'b0;
         RESULT_788 <= 16'b0;
         RESULT_789 <= 16'b0;
         RESULT_790 <= 16'b0;
         RESULT_791 <= 16'b0;
         RESULT_792 <= 16'b0;
         RESULT_793 <= 16'b0;
         RESULT_794 <= 16'b0;
         RESULT_795 <= 16'b0;
         RESULT_796 <= 16'b0;
         RESULT_797 <= 16'b0;
         RESULT_798 <= 16'b0;
         RESULT_799 <= 16'b0;
         RESULT_800 <= 16'b0;
         RESULT_801 <= 16'b0;
         RESULT_802 <= 16'b0;
         RESULT_803 <= 16'b0;
         RESULT_804 <= 16'b0;
         RESULT_805 <= 16'b0;
         RESULT_806 <= 16'b0;
         RESULT_807 <= 16'b0;
         RESULT_808 <= 16'b0;
         RESULT_809 <= 16'b0;
         RESULT_810 <= 16'b0;
         RESULT_811 <= 16'b0;
         RESULT_812 <= 16'b0;
         RESULT_813 <= 16'b0;
         RESULT_814 <= 16'b0;
         RESULT_815 <= 16'b0;
         RESULT_816 <= 16'b0;
         RESULT_817 <= 16'b0;
         RESULT_818 <= 16'b0;
         RESULT_819 <= 16'b0;
         RESULT_820 <= 16'b0;
         RESULT_821 <= 16'b0;
         RESULT_822 <= 16'b0;
         RESULT_823 <= 16'b0;
         RESULT_824 <= 16'b0;
         RESULT_825 <= 16'b0;
         RESULT_826 <= 16'b0;
         RESULT_827 <= 16'b0;
         RESULT_828 <= 16'b0;
         RESULT_829 <= 16'b0;
         RESULT_830 <= 16'b0;
         RESULT_831 <= 16'b0;
         RESULT_832 <= 16'b0;
         RESULT_833 <= 16'b0;
         RESULT_834 <= 16'b0;
         RESULT_835 <= 16'b0;
         RESULT_836 <= 16'b0;
         RESULT_837 <= 16'b0;
         RESULT_838 <= 16'b0;
         RESULT_839 <= 16'b0;
         RESULT_840 <= 16'b0;
         RESULT_841 <= 16'b0;
         RESULT_842 <= 16'b0;
         RESULT_843 <= 16'b0;
         RESULT_844 <= 16'b0;
         RESULT_845 <= 16'b0;
         RESULT_846 <= 16'b0;
         RESULT_847 <= 16'b0;
         RESULT_848 <= 16'b0;
         RESULT_849 <= 16'b0;
         RESULT_850 <= 16'b0;
         RESULT_851 <= 16'b0;
         RESULT_852 <= 16'b0;
         RESULT_853 <= 16'b0;
         RESULT_854 <= 16'b0;
         RESULT_855 <= 16'b0;
         RESULT_856 <= 16'b0;
         RESULT_857 <= 16'b0;
         RESULT_858 <= 16'b0;
         RESULT_859 <= 16'b0;
         RESULT_860 <= 16'b0;
         RESULT_861 <= 16'b0;
         RESULT_862 <= 16'b0;
         RESULT_863 <= 16'b0;
         RESULT_864 <= 16'b0;
         RESULT_865 <= 16'b0;
         RESULT_866 <= 16'b0;
         RESULT_867 <= 16'b0;
         RESULT_868 <= 16'b0;
         RESULT_869 <= 16'b0;
         RESULT_870 <= 16'b0;
         RESULT_871 <= 16'b0;
         RESULT_872 <= 16'b0;
         RESULT_873 <= 16'b0;
         RESULT_874 <= 16'b0;
         RESULT_875 <= 16'b0;
         RESULT_876 <= 16'b0;
         RESULT_877 <= 16'b0;
         RESULT_878 <= 16'b0;
         RESULT_879 <= 16'b0;
         RESULT_880 <= 16'b0;
         RESULT_881 <= 16'b0;
         RESULT_882 <= 16'b0;
         RESULT_883 <= 16'b0;
         RESULT_884 <= 16'b0;
         RESULT_885 <= 16'b0;
         RESULT_886 <= 16'b0;
         RESULT_887 <= 16'b0;
         RESULT_888 <= 16'b0;
         RESULT_889 <= 16'b0;
         RESULT_890 <= 16'b0;
         RESULT_891 <= 16'b0;
         RESULT_892 <= 16'b0;
         RESULT_893 <= 16'b0;
         RESULT_894 <= 16'b0;
         RESULT_895 <= 16'b0;
	  end
   end
   
   // Done signal and cycle counter
    always @(posedge CLK or negedge RSTN) begin
        if (!RSTN) begin
            count <= 0;
			case_enable <= 0;
        end else if (result_enable) begin
                if (count == 41) begin
					count <=0;
					case_enable <= 1;
                end else begin
                    count <= count + 1;
					case_enable <= 1;
                end
		end else begin
			count <= 0;
			case_enable <= 0;
		end
	end
         





endmodule

